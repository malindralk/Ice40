// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 15 2022 06:07:59

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    Y,
    mclock,
    DIGIT1,
    DIGIT2,
    DIGIT3,
    DIGIT4);

    output [7:0] Y;
    input mclock;
    output DIGIT1;
    output DIGIT2;
    output DIGIT3;
    output DIGIT4;

    wire N__2101;
    wire N__2100;
    wire N__2099;
    wire N__2090;
    wire N__2089;
    wire N__2088;
    wire N__2081;
    wire N__2080;
    wire N__2079;
    wire N__2072;
    wire N__2071;
    wire N__2070;
    wire N__2063;
    wire N__2062;
    wire N__2061;
    wire N__2054;
    wire N__2053;
    wire N__2052;
    wire N__2045;
    wire N__2044;
    wire N__2043;
    wire N__2036;
    wire N__2035;
    wire N__2034;
    wire N__2027;
    wire N__2026;
    wire N__2025;
    wire N__2018;
    wire N__2017;
    wire N__2016;
    wire N__2009;
    wire N__2008;
    wire N__2007;
    wire N__2000;
    wire N__1999;
    wire N__1998;
    wire N__1991;
    wire N__1990;
    wire N__1989;
    wire N__1972;
    wire N__1969;
    wire N__1966;
    wire N__1963;
    wire N__1960;
    wire N__1957;
    wire N__1954;
    wire N__1951;
    wire N__1948;
    wire N__1945;
    wire N__1942;
    wire N__1939;
    wire N__1936;
    wire N__1933;
    wire N__1930;
    wire N__1927;
    wire N__1924;
    wire N__1921;
    wire N__1920;
    wire N__1919;
    wire N__1918;
    wire N__1909;
    wire N__1908;
    wire N__1905;
    wire N__1904;
    wire N__1903;
    wire N__1902;
    wire N__1899;
    wire N__1898;
    wire N__1895;
    wire N__1892;
    wire N__1885;
    wire N__1882;
    wire N__1881;
    wire N__1880;
    wire N__1879;
    wire N__1872;
    wire N__1867;
    wire N__1864;
    wire N__1861;
    wire N__1852;
    wire N__1851;
    wire N__1848;
    wire N__1847;
    wire N__1846;
    wire N__1843;
    wire N__1834;
    wire N__1831;
    wire N__1830;
    wire N__1829;
    wire N__1828;
    wire N__1827;
    wire N__1824;
    wire N__1815;
    wire N__1814;
    wire N__1813;
    wire N__1812;
    wire N__1811;
    wire N__1808;
    wire N__1805;
    wire N__1800;
    wire N__1797;
    wire N__1794;
    wire N__1783;
    wire N__1782;
    wire N__1781;
    wire N__1780;
    wire N__1779;
    wire N__1778;
    wire N__1769;
    wire N__1768;
    wire N__1765;
    wire N__1762;
    wire N__1761;
    wire N__1758;
    wire N__1749;
    wire N__1748;
    wire N__1745;
    wire N__1742;
    wire N__1741;
    wire N__1740;
    wire N__1737;
    wire N__1734;
    wire N__1731;
    wire N__1728;
    wire N__1723;
    wire N__1714;
    wire N__1713;
    wire N__1710;
    wire N__1707;
    wire N__1706;
    wire N__1699;
    wire N__1696;
    wire N__1695;
    wire N__1694;
    wire N__1693;
    wire N__1692;
    wire N__1691;
    wire N__1688;
    wire N__1679;
    wire N__1678;
    wire N__1675;
    wire N__1674;
    wire N__1673;
    wire N__1670;
    wire N__1667;
    wire N__1664;
    wire N__1661;
    wire N__1656;
    wire N__1645;
    wire N__1642;
    wire N__1639;
    wire N__1636;
    wire N__1633;
    wire N__1630;
    wire N__1627;
    wire N__1624;
    wire N__1623;
    wire N__1620;
    wire N__1617;
    wire N__1612;
    wire N__1609;
    wire N__1608;
    wire N__1605;
    wire N__1602;
    wire N__1597;
    wire N__1596;
    wire N__1593;
    wire N__1590;
    wire N__1585;
    wire N__1584;
    wire N__1583;
    wire N__1582;
    wire N__1581;
    wire N__1580;
    wire N__1579;
    wire N__1578;
    wire N__1561;
    wire N__1558;
    wire N__1555;
    wire N__1552;
    wire N__1551;
    wire N__1550;
    wire N__1547;
    wire N__1544;
    wire N__1541;
    wire N__1538;
    wire N__1535;
    wire N__1532;
    wire N__1527;
    wire N__1522;
    wire N__1519;
    wire N__1516;
    wire N__1513;
    wire N__1510;
    wire N__1507;
    wire N__1506;
    wire N__1503;
    wire N__1500;
    wire N__1497;
    wire N__1492;
    wire N__1489;
    wire N__1488;
    wire N__1485;
    wire N__1482;
    wire N__1479;
    wire N__1474;
    wire N__1471;
    wire N__1470;
    wire N__1467;
    wire N__1464;
    wire N__1461;
    wire N__1456;
    wire N__1453;
    wire N__1452;
    wire N__1449;
    wire N__1446;
    wire N__1443;
    wire N__1438;
    wire N__1435;
    wire N__1434;
    wire N__1431;
    wire N__1428;
    wire N__1425;
    wire N__1420;
    wire N__1417;
    wire N__1416;
    wire N__1413;
    wire N__1410;
    wire N__1407;
    wire N__1402;
    wire N__1399;
    wire N__1398;
    wire N__1395;
    wire N__1392;
    wire N__1389;
    wire N__1384;
    wire N__1381;
    wire N__1380;
    wire N__1377;
    wire N__1374;
    wire N__1371;
    wire N__1366;
    wire N__1365;
    wire N__1362;
    wire N__1359;
    wire N__1356;
    wire N__1351;
    wire N__1348;
    wire N__1347;
    wire N__1344;
    wire N__1341;
    wire N__1338;
    wire N__1333;
    wire N__1330;
    wire N__1329;
    wire N__1326;
    wire N__1323;
    wire N__1320;
    wire N__1315;
    wire N__1312;
    wire N__1311;
    wire N__1308;
    wire N__1305;
    wire N__1302;
    wire N__1297;
    wire N__1294;
    wire N__1293;
    wire N__1290;
    wire N__1287;
    wire N__1284;
    wire N__1279;
    wire N__1278;
    wire N__1275;
    wire N__1272;
    wire N__1269;
    wire N__1264;
    wire N__1261;
    wire N__1260;
    wire N__1257;
    wire N__1254;
    wire N__1251;
    wire N__1246;
    wire N__1243;
    wire N__1242;
    wire N__1239;
    wire N__1236;
    wire N__1233;
    wire N__1228;
    wire N__1225;
    wire N__1224;
    wire N__1221;
    wire N__1218;
    wire N__1215;
    wire N__1210;
    wire N__1207;
    wire N__1204;
    wire N__1201;
    wire N__1200;
    wire N__1199;
    wire N__1196;
    wire N__1195;
    wire N__1190;
    wire N__1187;
    wire N__1184;
    wire N__1177;
    wire N__1176;
    wire N__1175;
    wire N__1172;
    wire N__1169;
    wire N__1166;
    wire N__1163;
    wire N__1160;
    wire N__1153;
    wire N__1150;
    wire N__1149;
    wire N__1146;
    wire N__1143;
    wire N__1140;
    wire N__1135;
    wire N__1134;
    wire N__1131;
    wire N__1128;
    wire N__1125;
    wire N__1120;
    wire N__1117;
    wire N__1116;
    wire N__1113;
    wire N__1110;
    wire N__1107;
    wire N__1102;
    wire N__1099;
    wire N__1098;
    wire N__1095;
    wire N__1092;
    wire N__1089;
    wire N__1084;
    wire N__1081;
    wire N__1080;
    wire N__1077;
    wire N__1074;
    wire N__1071;
    wire N__1066;
    wire N__1063;
    wire N__1062;
    wire N__1059;
    wire N__1056;
    wire N__1053;
    wire N__1048;
    wire N__1045;
    wire N__1042;
    wire N__1039;
    wire N__1036;
    wire N__1033;
    wire N__1030;
    wire N__1027;
    wire N__1024;
    wire N__1021;
    wire N__1018;
    wire N__1015;
    wire N__1012;
    wire N__1009;
    wire N__1006;
    wire N__1003;
    wire N__1000;
    wire N__997;
    wire N__994;
    wire N__991;
    wire N__988;
    wire GNDG0;
    wire VCCG0;
    wire bfn_22_17_0_;
    wire un2_cntdiv_cry_1;
    wire un2_cntdiv_cry_2;
    wire un2_cntdiv_cry_3;
    wire un2_cntdiv_cry_4;
    wire un2_cntdiv_cry_5;
    wire un2_cntdiv_cry_6;
    wire un2_cntdiv_cry_7;
    wire un2_cntdiv_cry_8;
    wire bfn_22_18_0_;
    wire un2_cntdiv_cry_9;
    wire un2_cntdiv_cry_10;
    wire un2_cntdiv_cry_11;
    wire un2_cntdiv_cry_12;
    wire un2_cntdiv_cry_13;
    wire un2_cntdiv_cry_14;
    wire un2_cntdiv_cry_15;
    wire un2_cntdiv_cry_16;
    wire bfn_22_19_0_;
    wire un2_cntdiv_cry_17;
    wire un2_cntdiv_cry_18;
    wire un2_cntdiv_cry_19;
    wire un2_cntdiv_cry_20;
    wire un2_cntdiv_cry_21;
    wire un2_cntdiv_cry_22;
    wire un2_cntdiv_cry_23;
    wire cntDivZ0Z_0;
    wire cntDivZ0Z_1;
    wire bfn_22_20_0_;
    wire cntDivZ0Z_2;
    wire un2_cntdiv_1_cry_1;
    wire cntDivZ0Z_3;
    wire un2_cntdiv_1_cry_2;
    wire cntDivZ0Z_4;
    wire un2_cntdiv_1_cry_3;
    wire cntDivZ0Z_5;
    wire un2_cntdiv_1_cry_4;
    wire cntDivZ0Z_6;
    wire un2_cntdiv_1_cry_5;
    wire cntDivZ0Z_7;
    wire un2_cntdiv_1_cry_6;
    wire cntDivZ0Z_8;
    wire un2_cntdiv_1_cry_7;
    wire un2_cntdiv_1_cry_8;
    wire cntDivZ0Z_9;
    wire bfn_22_21_0_;
    wire cntDivZ0Z_10;
    wire un2_cntdiv_1_cry_9;
    wire cntDivZ0Z_11;
    wire un2_cntdiv_1_cry_10;
    wire cntDivZ0Z_12;
    wire un2_cntdiv_1_cry_11;
    wire cntDivZ0Z_13;
    wire un2_cntdiv_1_cry_12;
    wire cntDivZ0Z_14;
    wire un2_cntdiv_1_cry_13;
    wire cntDivZ0Z_15;
    wire un2_cntdiv_1_cry_14;
    wire cntDivZ0Z_16;
    wire un2_cntdiv_1_cry_15;
    wire un2_cntdiv_1_cry_16;
    wire cntDivZ0Z_17;
    wire bfn_22_22_0_;
    wire cntDivZ0Z_18;
    wire un2_cntdiv_1_cry_17;
    wire cntDivZ0Z_19;
    wire un2_cntdiv_1_cry_18;
    wire cntDivZ0Z_20;
    wire un2_cntdiv_1_cry_19;
    wire cntDivZ0Z_21;
    wire un2_cntdiv_1_cry_20;
    wire cntDivZ0Z_22;
    wire un2_cntdiv_1_cry_21;
    wire cntDivZ0Z_23;
    wire un2_cntdiv_1_cry_22;
    wire cntDivZ0Z_24;
    wire un2_cntdiv_1_cry_23;
    wire un2_cntdiv_1_cry_24;
    wire bfn_22_23_0_;
    wire un2_cntdiv_1_cry_24_c_RNI73PBZ0;
    wire cntDiv_i_25;
    wire mclock_0_c_g;
    wire cntDiv_RNIETOHZ0Z_25;
    wire Y_c_1;
    wire Y_c_4;
    wire Y_c_0;
    wire Y_c_2;
    wire Y_c_7;
    wire Y_c_6;
    wire Y_c_3;
    wire value_1;
    wire value_3;
    wire value_2;
    wire value_0;
    wire Y_c_5;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    PRE_IO_GBUF mclock_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2099),
            .GLOBALBUFFEROUTPUT(mclock_0_c_g));
    IO_PAD mclock_ibuf_gb_io_iopad (
            .OE(N__2101),
            .DIN(N__2100),
            .DOUT(N__2099),
            .PACKAGEPIN(mclock));
    defparam mclock_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam mclock_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO mclock_ibuf_gb_io_preio (
            .PADOEN(N__2101),
            .PADOUT(N__2100),
            .PADIN(N__2099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_7_iopad (
            .OE(N__2090),
            .DIN(N__2089),
            .DOUT(N__2088),
            .PACKAGEPIN(Y[7]));
    defparam Y_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_7_preio (
            .PADOEN(N__2090),
            .PADOUT(N__2089),
            .PADIN(N__2088),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1948),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_0_iopad (
            .OE(N__2081),
            .DIN(N__2080),
            .DOUT(N__2079),
            .PACKAGEPIN(Y[0]));
    defparam Y_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_0_preio (
            .PADOEN(N__2081),
            .PADOUT(N__2080),
            .PADIN(N__2079),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1972),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DIGIT2_obuf_iopad (
            .OE(N__2072),
            .DIN(N__2071),
            .DOUT(N__2070),
            .PACKAGEPIN(DIGIT2));
    defparam DIGIT2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DIGIT2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DIGIT2_obuf_preio (
            .PADOEN(N__2072),
            .PADOUT(N__2071),
            .PADIN(N__2070),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_4_iopad (
            .OE(N__2063),
            .DIN(N__2062),
            .DOUT(N__2061),
            .PACKAGEPIN(Y[4]));
    defparam Y_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_4_preio (
            .PADOEN(N__2063),
            .PADOUT(N__2062),
            .PADIN(N__2061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1516),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DIGIT1_obuf_iopad (
            .OE(N__2054),
            .DIN(N__2053),
            .DOUT(N__2052),
            .PACKAGEPIN(DIGIT1));
    defparam DIGIT1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DIGIT1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DIGIT1_obuf_preio (
            .PADOEN(N__2054),
            .PADOUT(N__2053),
            .PADIN(N__2052),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1633),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_1_iopad (
            .OE(N__2045),
            .DIN(N__2044),
            .DOUT(N__2043),
            .PACKAGEPIN(Y[1]));
    defparam Y_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_1_preio (
            .PADOEN(N__2045),
            .PADOUT(N__2044),
            .PADIN(N__2043),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1522),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_5_iopad (
            .OE(N__2036),
            .DIN(N__2035),
            .DOUT(N__2034),
            .PACKAGEPIN(Y[5]));
    defparam Y_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_5_preio (
            .PADOEN(N__2036),
            .PADOUT(N__2035),
            .PADIN(N__2034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1645),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DIGIT3_obuf_iopad (
            .OE(N__2027),
            .DIN(N__2026),
            .DOUT(N__2025),
            .PACKAGEPIN(DIGIT3));
    defparam DIGIT3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DIGIT3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DIGIT3_obuf_preio (
            .PADOEN(N__2027),
            .PADOUT(N__2026),
            .PADIN(N__2025),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1623),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_2_iopad (
            .OE(N__2018),
            .DIN(N__2017),
            .DOUT(N__2016),
            .PACKAGEPIN(Y[2]));
    defparam Y_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_2_preio (
            .PADOEN(N__2018),
            .PADOUT(N__2017),
            .PADIN(N__2016),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1960),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DIGIT4_obuf_iopad (
            .OE(N__2009),
            .DIN(N__2008),
            .DOUT(N__2007),
            .PACKAGEPIN(DIGIT4));
    defparam DIGIT4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DIGIT4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DIGIT4_obuf_preio (
            .PADOEN(N__2009),
            .PADOUT(N__2008),
            .PADIN(N__2007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_6_iopad (
            .OE(N__2000),
            .DIN(N__1999),
            .DOUT(N__1998),
            .PACKAGEPIN(Y[6]));
    defparam Y_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_6_preio (
            .PADOEN(N__2000),
            .PADOUT(N__1999),
            .PADIN(N__1998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD Y_obuf_3_iopad (
            .OE(N__1991),
            .DIN(N__1990),
            .DOUT(N__1989),
            .PACKAGEPIN(Y[3]));
    defparam Y_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam Y_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO Y_obuf_3_preio (
            .PADOEN(N__1991),
            .PADOUT(N__1990),
            .PADIN(N__1989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1927),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__417 (
            .O(N__1972),
            .I(N__1969));
    LocalMux I__416 (
            .O(N__1969),
            .I(N__1966));
    Span4Mux_s0_h I__415 (
            .O(N__1966),
            .I(N__1963));
    Odrv4 I__414 (
            .O(N__1963),
            .I(Y_c_0));
    IoInMux I__413 (
            .O(N__1960),
            .I(N__1957));
    LocalMux I__412 (
            .O(N__1957),
            .I(N__1954));
    Span4Mux_s0_h I__411 (
            .O(N__1954),
            .I(N__1951));
    Odrv4 I__410 (
            .O(N__1951),
            .I(Y_c_2));
    IoInMux I__409 (
            .O(N__1948),
            .I(N__1945));
    LocalMux I__408 (
            .O(N__1945),
            .I(N__1942));
    Span4Mux_s1_h I__407 (
            .O(N__1942),
            .I(N__1939));
    Span4Mux_v I__406 (
            .O(N__1939),
            .I(N__1936));
    Odrv4 I__405 (
            .O(N__1936),
            .I(Y_c_7));
    IoInMux I__404 (
            .O(N__1933),
            .I(N__1930));
    LocalMux I__403 (
            .O(N__1930),
            .I(Y_c_6));
    IoInMux I__402 (
            .O(N__1927),
            .I(N__1924));
    LocalMux I__401 (
            .O(N__1924),
            .I(Y_c_3));
    InMux I__400 (
            .O(N__1921),
            .I(N__1909));
    InMux I__399 (
            .O(N__1920),
            .I(N__1909));
    InMux I__398 (
            .O(N__1919),
            .I(N__1909));
    InMux I__397 (
            .O(N__1918),
            .I(N__1909));
    LocalMux I__396 (
            .O(N__1909),
            .I(N__1905));
    CascadeMux I__395 (
            .O(N__1908),
            .I(N__1899));
    Span4Mux_v I__394 (
            .O(N__1905),
            .I(N__1895));
    InMux I__393 (
            .O(N__1904),
            .I(N__1892));
    InMux I__392 (
            .O(N__1903),
            .I(N__1885));
    InMux I__391 (
            .O(N__1902),
            .I(N__1885));
    InMux I__390 (
            .O(N__1899),
            .I(N__1885));
    CascadeMux I__389 (
            .O(N__1898),
            .I(N__1882));
    Sp12to4 I__388 (
            .O(N__1895),
            .I(N__1872));
    LocalMux I__387 (
            .O(N__1892),
            .I(N__1872));
    LocalMux I__386 (
            .O(N__1885),
            .I(N__1872));
    InMux I__385 (
            .O(N__1882),
            .I(N__1867));
    InMux I__384 (
            .O(N__1881),
            .I(N__1867));
    InMux I__383 (
            .O(N__1880),
            .I(N__1864));
    InMux I__382 (
            .O(N__1879),
            .I(N__1861));
    Odrv12 I__381 (
            .O(N__1872),
            .I(value_1));
    LocalMux I__380 (
            .O(N__1867),
            .I(value_1));
    LocalMux I__379 (
            .O(N__1864),
            .I(value_1));
    LocalMux I__378 (
            .O(N__1861),
            .I(value_1));
    CascadeMux I__377 (
            .O(N__1852),
            .I(N__1848));
    CascadeMux I__376 (
            .O(N__1851),
            .I(N__1843));
    InMux I__375 (
            .O(N__1848),
            .I(N__1834));
    InMux I__374 (
            .O(N__1847),
            .I(N__1834));
    InMux I__373 (
            .O(N__1846),
            .I(N__1834));
    InMux I__372 (
            .O(N__1843),
            .I(N__1834));
    LocalMux I__371 (
            .O(N__1834),
            .I(N__1831));
    Span4Mux_v I__370 (
            .O(N__1831),
            .I(N__1824));
    InMux I__369 (
            .O(N__1830),
            .I(N__1815));
    InMux I__368 (
            .O(N__1829),
            .I(N__1815));
    InMux I__367 (
            .O(N__1828),
            .I(N__1815));
    InMux I__366 (
            .O(N__1827),
            .I(N__1815));
    Span4Mux_h I__365 (
            .O(N__1824),
            .I(N__1808));
    LocalMux I__364 (
            .O(N__1815),
            .I(N__1805));
    InMux I__363 (
            .O(N__1814),
            .I(N__1800));
    InMux I__362 (
            .O(N__1813),
            .I(N__1800));
    InMux I__361 (
            .O(N__1812),
            .I(N__1797));
    InMux I__360 (
            .O(N__1811),
            .I(N__1794));
    Odrv4 I__359 (
            .O(N__1808),
            .I(value_3));
    Odrv12 I__358 (
            .O(N__1805),
            .I(value_3));
    LocalMux I__357 (
            .O(N__1800),
            .I(value_3));
    LocalMux I__356 (
            .O(N__1797),
            .I(value_3));
    LocalMux I__355 (
            .O(N__1794),
            .I(value_3));
    InMux I__354 (
            .O(N__1783),
            .I(N__1769));
    InMux I__353 (
            .O(N__1782),
            .I(N__1769));
    InMux I__352 (
            .O(N__1781),
            .I(N__1769));
    InMux I__351 (
            .O(N__1780),
            .I(N__1769));
    CascadeMux I__350 (
            .O(N__1779),
            .I(N__1765));
    CascadeMux I__349 (
            .O(N__1778),
            .I(N__1762));
    LocalMux I__348 (
            .O(N__1769),
            .I(N__1758));
    InMux I__347 (
            .O(N__1768),
            .I(N__1749));
    InMux I__346 (
            .O(N__1765),
            .I(N__1749));
    InMux I__345 (
            .O(N__1762),
            .I(N__1749));
    InMux I__344 (
            .O(N__1761),
            .I(N__1749));
    Span4Mux_v I__343 (
            .O(N__1758),
            .I(N__1745));
    LocalMux I__342 (
            .O(N__1749),
            .I(N__1742));
    CascadeMux I__341 (
            .O(N__1748),
            .I(N__1737));
    Span4Mux_h I__340 (
            .O(N__1745),
            .I(N__1734));
    Span12Mux_s2_h I__339 (
            .O(N__1742),
            .I(N__1731));
    InMux I__338 (
            .O(N__1741),
            .I(N__1728));
    InMux I__337 (
            .O(N__1740),
            .I(N__1723));
    InMux I__336 (
            .O(N__1737),
            .I(N__1723));
    Odrv4 I__335 (
            .O(N__1734),
            .I(value_2));
    Odrv12 I__334 (
            .O(N__1731),
            .I(value_2));
    LocalMux I__333 (
            .O(N__1728),
            .I(value_2));
    LocalMux I__332 (
            .O(N__1723),
            .I(value_2));
    CascadeMux I__331 (
            .O(N__1714),
            .I(N__1710));
    CascadeMux I__330 (
            .O(N__1713),
            .I(N__1707));
    InMux I__329 (
            .O(N__1710),
            .I(N__1699));
    InMux I__328 (
            .O(N__1707),
            .I(N__1699));
    InMux I__327 (
            .O(N__1706),
            .I(N__1699));
    LocalMux I__326 (
            .O(N__1699),
            .I(N__1696));
    Span4Mux_s3_h I__325 (
            .O(N__1696),
            .I(N__1688));
    InMux I__324 (
            .O(N__1695),
            .I(N__1679));
    InMux I__323 (
            .O(N__1694),
            .I(N__1679));
    InMux I__322 (
            .O(N__1693),
            .I(N__1679));
    InMux I__321 (
            .O(N__1692),
            .I(N__1679));
    CascadeMux I__320 (
            .O(N__1691),
            .I(N__1675));
    Span4Mux_h I__319 (
            .O(N__1688),
            .I(N__1670));
    LocalMux I__318 (
            .O(N__1679),
            .I(N__1667));
    InMux I__317 (
            .O(N__1678),
            .I(N__1664));
    InMux I__316 (
            .O(N__1675),
            .I(N__1661));
    InMux I__315 (
            .O(N__1674),
            .I(N__1656));
    InMux I__314 (
            .O(N__1673),
            .I(N__1656));
    Odrv4 I__313 (
            .O(N__1670),
            .I(value_0));
    Odrv12 I__312 (
            .O(N__1667),
            .I(value_0));
    LocalMux I__311 (
            .O(N__1664),
            .I(value_0));
    LocalMux I__310 (
            .O(N__1661),
            .I(value_0));
    LocalMux I__309 (
            .O(N__1656),
            .I(value_0));
    IoInMux I__308 (
            .O(N__1645),
            .I(N__1642));
    LocalMux I__307 (
            .O(N__1642),
            .I(N__1639));
    Span12Mux_s0_h I__306 (
            .O(N__1639),
            .I(N__1636));
    Odrv12 I__305 (
            .O(N__1636),
            .I(Y_c_5));
    IoInMux I__304 (
            .O(N__1633),
            .I(N__1630));
    LocalMux I__303 (
            .O(N__1630),
            .I(N__1627));
    IoSpan4Mux I__302 (
            .O(N__1627),
            .I(N__1624));
    Span4Mux_s2_v I__301 (
            .O(N__1624),
            .I(N__1620));
    IoInMux I__300 (
            .O(N__1623),
            .I(N__1617));
    Odrv4 I__299 (
            .O(N__1620),
            .I(CONSTANT_ONE_NET));
    LocalMux I__298 (
            .O(N__1617),
            .I(CONSTANT_ONE_NET));
    InMux I__297 (
            .O(N__1612),
            .I(bfn_22_23_0_));
    InMux I__296 (
            .O(N__1609),
            .I(N__1605));
    InMux I__295 (
            .O(N__1608),
            .I(N__1602));
    LocalMux I__294 (
            .O(N__1605),
            .I(un2_cntdiv_1_cry_24_c_RNI73PBZ0));
    LocalMux I__293 (
            .O(N__1602),
            .I(un2_cntdiv_1_cry_24_c_RNI73PBZ0));
    InMux I__292 (
            .O(N__1597),
            .I(N__1593));
    InMux I__291 (
            .O(N__1596),
            .I(N__1590));
    LocalMux I__290 (
            .O(N__1593),
            .I(cntDiv_i_25));
    LocalMux I__289 (
            .O(N__1590),
            .I(cntDiv_i_25));
    ClkMux I__288 (
            .O(N__1585),
            .I(N__1561));
    ClkMux I__287 (
            .O(N__1584),
            .I(N__1561));
    ClkMux I__286 (
            .O(N__1583),
            .I(N__1561));
    ClkMux I__285 (
            .O(N__1582),
            .I(N__1561));
    ClkMux I__284 (
            .O(N__1581),
            .I(N__1561));
    ClkMux I__283 (
            .O(N__1580),
            .I(N__1561));
    ClkMux I__282 (
            .O(N__1579),
            .I(N__1561));
    ClkMux I__281 (
            .O(N__1578),
            .I(N__1561));
    GlobalMux I__280 (
            .O(N__1561),
            .I(N__1558));
    gio2CtrlBuf I__279 (
            .O(N__1558),
            .I(mclock_0_c_g));
    CEMux I__278 (
            .O(N__1555),
            .I(N__1552));
    LocalMux I__277 (
            .O(N__1552),
            .I(N__1547));
    CEMux I__276 (
            .O(N__1551),
            .I(N__1544));
    CEMux I__275 (
            .O(N__1550),
            .I(N__1541));
    Span4Mux_h I__274 (
            .O(N__1547),
            .I(N__1538));
    LocalMux I__273 (
            .O(N__1544),
            .I(N__1535));
    LocalMux I__272 (
            .O(N__1541),
            .I(N__1532));
    Span4Mux_h I__271 (
            .O(N__1538),
            .I(N__1527));
    Span4Mux_h I__270 (
            .O(N__1535),
            .I(N__1527));
    Odrv12 I__269 (
            .O(N__1532),
            .I(cntDiv_RNIETOHZ0Z_25));
    Odrv4 I__268 (
            .O(N__1527),
            .I(cntDiv_RNIETOHZ0Z_25));
    IoInMux I__267 (
            .O(N__1522),
            .I(N__1519));
    LocalMux I__266 (
            .O(N__1519),
            .I(Y_c_1));
    IoInMux I__265 (
            .O(N__1516),
            .I(N__1513));
    LocalMux I__264 (
            .O(N__1513),
            .I(Y_c_4));
    CascadeMux I__263 (
            .O(N__1510),
            .I(N__1507));
    InMux I__262 (
            .O(N__1507),
            .I(N__1503));
    InMux I__261 (
            .O(N__1506),
            .I(N__1500));
    LocalMux I__260 (
            .O(N__1503),
            .I(N__1497));
    LocalMux I__259 (
            .O(N__1500),
            .I(cntDivZ0Z_16));
    Odrv4 I__258 (
            .O(N__1497),
            .I(cntDivZ0Z_16));
    CascadeMux I__257 (
            .O(N__1492),
            .I(N__1489));
    InMux I__256 (
            .O(N__1489),
            .I(N__1485));
    InMux I__255 (
            .O(N__1488),
            .I(N__1482));
    LocalMux I__254 (
            .O(N__1485),
            .I(N__1479));
    LocalMux I__253 (
            .O(N__1482),
            .I(cntDivZ0Z_17));
    Odrv12 I__252 (
            .O(N__1479),
            .I(cntDivZ0Z_17));
    CascadeMux I__251 (
            .O(N__1474),
            .I(N__1471));
    InMux I__250 (
            .O(N__1471),
            .I(N__1467));
    InMux I__249 (
            .O(N__1470),
            .I(N__1464));
    LocalMux I__248 (
            .O(N__1467),
            .I(N__1461));
    LocalMux I__247 (
            .O(N__1464),
            .I(cntDivZ0Z_18));
    Odrv12 I__246 (
            .O(N__1461),
            .I(cntDivZ0Z_18));
    CascadeMux I__245 (
            .O(N__1456),
            .I(N__1453));
    InMux I__244 (
            .O(N__1453),
            .I(N__1449));
    InMux I__243 (
            .O(N__1452),
            .I(N__1446));
    LocalMux I__242 (
            .O(N__1449),
            .I(N__1443));
    LocalMux I__241 (
            .O(N__1446),
            .I(cntDivZ0Z_19));
    Odrv4 I__240 (
            .O(N__1443),
            .I(cntDivZ0Z_19));
    CascadeMux I__239 (
            .O(N__1438),
            .I(N__1435));
    InMux I__238 (
            .O(N__1435),
            .I(N__1431));
    InMux I__237 (
            .O(N__1434),
            .I(N__1428));
    LocalMux I__236 (
            .O(N__1431),
            .I(N__1425));
    LocalMux I__235 (
            .O(N__1428),
            .I(cntDivZ0Z_20));
    Odrv4 I__234 (
            .O(N__1425),
            .I(cntDivZ0Z_20));
    CascadeMux I__233 (
            .O(N__1420),
            .I(N__1417));
    InMux I__232 (
            .O(N__1417),
            .I(N__1413));
    InMux I__231 (
            .O(N__1416),
            .I(N__1410));
    LocalMux I__230 (
            .O(N__1413),
            .I(N__1407));
    LocalMux I__229 (
            .O(N__1410),
            .I(cntDivZ0Z_21));
    Odrv4 I__228 (
            .O(N__1407),
            .I(cntDivZ0Z_21));
    CascadeMux I__227 (
            .O(N__1402),
            .I(N__1399));
    InMux I__226 (
            .O(N__1399),
            .I(N__1395));
    InMux I__225 (
            .O(N__1398),
            .I(N__1392));
    LocalMux I__224 (
            .O(N__1395),
            .I(N__1389));
    LocalMux I__223 (
            .O(N__1392),
            .I(cntDivZ0Z_22));
    Odrv4 I__222 (
            .O(N__1389),
            .I(cntDivZ0Z_22));
    CascadeMux I__221 (
            .O(N__1384),
            .I(N__1381));
    InMux I__220 (
            .O(N__1381),
            .I(N__1377));
    InMux I__219 (
            .O(N__1380),
            .I(N__1374));
    LocalMux I__218 (
            .O(N__1377),
            .I(N__1371));
    LocalMux I__217 (
            .O(N__1374),
            .I(cntDivZ0Z_23));
    Odrv4 I__216 (
            .O(N__1371),
            .I(cntDivZ0Z_23));
    InMux I__215 (
            .O(N__1366),
            .I(N__1362));
    InMux I__214 (
            .O(N__1365),
            .I(N__1359));
    LocalMux I__213 (
            .O(N__1362),
            .I(N__1356));
    LocalMux I__212 (
            .O(N__1359),
            .I(cntDivZ0Z_24));
    Odrv4 I__211 (
            .O(N__1356),
            .I(cntDivZ0Z_24));
    CascadeMux I__210 (
            .O(N__1351),
            .I(N__1348));
    InMux I__209 (
            .O(N__1348),
            .I(N__1344));
    InMux I__208 (
            .O(N__1347),
            .I(N__1341));
    LocalMux I__207 (
            .O(N__1344),
            .I(N__1338));
    LocalMux I__206 (
            .O(N__1341),
            .I(cntDivZ0Z_8));
    Odrv4 I__205 (
            .O(N__1338),
            .I(cntDivZ0Z_8));
    CascadeMux I__204 (
            .O(N__1333),
            .I(N__1330));
    InMux I__203 (
            .O(N__1330),
            .I(N__1326));
    InMux I__202 (
            .O(N__1329),
            .I(N__1323));
    LocalMux I__201 (
            .O(N__1326),
            .I(N__1320));
    LocalMux I__200 (
            .O(N__1323),
            .I(cntDivZ0Z_9));
    Odrv12 I__199 (
            .O(N__1320),
            .I(cntDivZ0Z_9));
    CascadeMux I__198 (
            .O(N__1315),
            .I(N__1312));
    InMux I__197 (
            .O(N__1312),
            .I(N__1308));
    InMux I__196 (
            .O(N__1311),
            .I(N__1305));
    LocalMux I__195 (
            .O(N__1308),
            .I(N__1302));
    LocalMux I__194 (
            .O(N__1305),
            .I(cntDivZ0Z_10));
    Odrv12 I__193 (
            .O(N__1302),
            .I(cntDivZ0Z_10));
    CascadeMux I__192 (
            .O(N__1297),
            .I(N__1294));
    InMux I__191 (
            .O(N__1294),
            .I(N__1290));
    InMux I__190 (
            .O(N__1293),
            .I(N__1287));
    LocalMux I__189 (
            .O(N__1290),
            .I(N__1284));
    LocalMux I__188 (
            .O(N__1287),
            .I(cntDivZ0Z_11));
    Odrv4 I__187 (
            .O(N__1284),
            .I(cntDivZ0Z_11));
    InMux I__186 (
            .O(N__1279),
            .I(N__1275));
    InMux I__185 (
            .O(N__1278),
            .I(N__1272));
    LocalMux I__184 (
            .O(N__1275),
            .I(N__1269));
    LocalMux I__183 (
            .O(N__1272),
            .I(cntDivZ0Z_12));
    Odrv4 I__182 (
            .O(N__1269),
            .I(cntDivZ0Z_12));
    CascadeMux I__181 (
            .O(N__1264),
            .I(N__1261));
    InMux I__180 (
            .O(N__1261),
            .I(N__1257));
    InMux I__179 (
            .O(N__1260),
            .I(N__1254));
    LocalMux I__178 (
            .O(N__1257),
            .I(N__1251));
    LocalMux I__177 (
            .O(N__1254),
            .I(cntDivZ0Z_13));
    Odrv4 I__176 (
            .O(N__1251),
            .I(cntDivZ0Z_13));
    CascadeMux I__175 (
            .O(N__1246),
            .I(N__1243));
    InMux I__174 (
            .O(N__1243),
            .I(N__1239));
    InMux I__173 (
            .O(N__1242),
            .I(N__1236));
    LocalMux I__172 (
            .O(N__1239),
            .I(N__1233));
    LocalMux I__171 (
            .O(N__1236),
            .I(cntDivZ0Z_14));
    Odrv4 I__170 (
            .O(N__1233),
            .I(cntDivZ0Z_14));
    CascadeMux I__169 (
            .O(N__1228),
            .I(N__1225));
    InMux I__168 (
            .O(N__1225),
            .I(N__1221));
    InMux I__167 (
            .O(N__1224),
            .I(N__1218));
    LocalMux I__166 (
            .O(N__1221),
            .I(N__1215));
    LocalMux I__165 (
            .O(N__1218),
            .I(cntDivZ0Z_15));
    Odrv4 I__164 (
            .O(N__1215),
            .I(cntDivZ0Z_15));
    InMux I__163 (
            .O(N__1210),
            .I(un2_cntdiv_cry_22));
    InMux I__162 (
            .O(N__1207),
            .I(un2_cntdiv_cry_23));
    CascadeMux I__161 (
            .O(N__1204),
            .I(N__1201));
    InMux I__160 (
            .O(N__1201),
            .I(N__1196));
    InMux I__159 (
            .O(N__1200),
            .I(N__1190));
    InMux I__158 (
            .O(N__1199),
            .I(N__1190));
    LocalMux I__157 (
            .O(N__1196),
            .I(N__1187));
    InMux I__156 (
            .O(N__1195),
            .I(N__1184));
    LocalMux I__155 (
            .O(N__1190),
            .I(cntDivZ0Z_0));
    Odrv4 I__154 (
            .O(N__1187),
            .I(cntDivZ0Z_0));
    LocalMux I__153 (
            .O(N__1184),
            .I(cntDivZ0Z_0));
    InMux I__152 (
            .O(N__1177),
            .I(N__1172));
    CascadeMux I__151 (
            .O(N__1176),
            .I(N__1169));
    InMux I__150 (
            .O(N__1175),
            .I(N__1166));
    LocalMux I__149 (
            .O(N__1172),
            .I(N__1163));
    InMux I__148 (
            .O(N__1169),
            .I(N__1160));
    LocalMux I__147 (
            .O(N__1166),
            .I(cntDivZ0Z_1));
    Odrv4 I__146 (
            .O(N__1163),
            .I(cntDivZ0Z_1));
    LocalMux I__145 (
            .O(N__1160),
            .I(cntDivZ0Z_1));
    CascadeMux I__144 (
            .O(N__1153),
            .I(N__1150));
    InMux I__143 (
            .O(N__1150),
            .I(N__1146));
    InMux I__142 (
            .O(N__1149),
            .I(N__1143));
    LocalMux I__141 (
            .O(N__1146),
            .I(N__1140));
    LocalMux I__140 (
            .O(N__1143),
            .I(cntDivZ0Z_2));
    Odrv12 I__139 (
            .O(N__1140),
            .I(cntDivZ0Z_2));
    InMux I__138 (
            .O(N__1135),
            .I(N__1131));
    InMux I__137 (
            .O(N__1134),
            .I(N__1128));
    LocalMux I__136 (
            .O(N__1131),
            .I(N__1125));
    LocalMux I__135 (
            .O(N__1128),
            .I(cntDivZ0Z_3));
    Odrv4 I__134 (
            .O(N__1125),
            .I(cntDivZ0Z_3));
    CascadeMux I__133 (
            .O(N__1120),
            .I(N__1117));
    InMux I__132 (
            .O(N__1117),
            .I(N__1113));
    InMux I__131 (
            .O(N__1116),
            .I(N__1110));
    LocalMux I__130 (
            .O(N__1113),
            .I(N__1107));
    LocalMux I__129 (
            .O(N__1110),
            .I(cntDivZ0Z_4));
    Odrv4 I__128 (
            .O(N__1107),
            .I(cntDivZ0Z_4));
    CascadeMux I__127 (
            .O(N__1102),
            .I(N__1099));
    InMux I__126 (
            .O(N__1099),
            .I(N__1095));
    InMux I__125 (
            .O(N__1098),
            .I(N__1092));
    LocalMux I__124 (
            .O(N__1095),
            .I(N__1089));
    LocalMux I__123 (
            .O(N__1092),
            .I(cntDivZ0Z_5));
    Odrv4 I__122 (
            .O(N__1089),
            .I(cntDivZ0Z_5));
    CascadeMux I__121 (
            .O(N__1084),
            .I(N__1081));
    InMux I__120 (
            .O(N__1081),
            .I(N__1077));
    InMux I__119 (
            .O(N__1080),
            .I(N__1074));
    LocalMux I__118 (
            .O(N__1077),
            .I(N__1071));
    LocalMux I__117 (
            .O(N__1074),
            .I(cntDivZ0Z_6));
    Odrv4 I__116 (
            .O(N__1071),
            .I(cntDivZ0Z_6));
    CascadeMux I__115 (
            .O(N__1066),
            .I(N__1063));
    InMux I__114 (
            .O(N__1063),
            .I(N__1059));
    InMux I__113 (
            .O(N__1062),
            .I(N__1056));
    LocalMux I__112 (
            .O(N__1059),
            .I(N__1053));
    LocalMux I__111 (
            .O(N__1056),
            .I(cntDivZ0Z_7));
    Odrv4 I__110 (
            .O(N__1053),
            .I(cntDivZ0Z_7));
    InMux I__109 (
            .O(N__1048),
            .I(un2_cntdiv_cry_13));
    InMux I__108 (
            .O(N__1045),
            .I(un2_cntdiv_cry_14));
    InMux I__107 (
            .O(N__1042),
            .I(un2_cntdiv_cry_15));
    InMux I__106 (
            .O(N__1039),
            .I(bfn_22_19_0_));
    InMux I__105 (
            .O(N__1036),
            .I(un2_cntdiv_cry_17));
    InMux I__104 (
            .O(N__1033),
            .I(un2_cntdiv_cry_18));
    InMux I__103 (
            .O(N__1030),
            .I(un2_cntdiv_cry_19));
    InMux I__102 (
            .O(N__1027),
            .I(un2_cntdiv_cry_20));
    InMux I__101 (
            .O(N__1024),
            .I(un2_cntdiv_cry_21));
    InMux I__100 (
            .O(N__1021),
            .I(un2_cntdiv_cry_4));
    InMux I__99 (
            .O(N__1018),
            .I(un2_cntdiv_cry_5));
    InMux I__98 (
            .O(N__1015),
            .I(un2_cntdiv_cry_6));
    InMux I__97 (
            .O(N__1012),
            .I(un2_cntdiv_cry_7));
    InMux I__96 (
            .O(N__1009),
            .I(bfn_22_18_0_));
    InMux I__95 (
            .O(N__1006),
            .I(un2_cntdiv_cry_9));
    InMux I__94 (
            .O(N__1003),
            .I(un2_cntdiv_cry_10));
    InMux I__93 (
            .O(N__1000),
            .I(un2_cntdiv_cry_11));
    InMux I__92 (
            .O(N__997),
            .I(un2_cntdiv_cry_12));
    InMux I__91 (
            .O(N__994),
            .I(un2_cntdiv_cry_1));
    InMux I__90 (
            .O(N__991),
            .I(un2_cntdiv_cry_2));
    InMux I__89 (
            .O(N__988),
            .I(un2_cntdiv_cry_3));
    defparam IN_MUX_bfv_22_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_17_0_));
    defparam IN_MUX_bfv_22_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_18_0_ (
            .carryinitin(un2_cntdiv_cry_8),
            .carryinitout(bfn_22_18_0_));
    defparam IN_MUX_bfv_22_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_19_0_ (
            .carryinitin(un2_cntdiv_cry_16),
            .carryinitout(bfn_22_19_0_));
    defparam IN_MUX_bfv_22_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_20_0_));
    defparam IN_MUX_bfv_22_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_21_0_ (
            .carryinitin(un2_cntdiv_1_cry_8),
            .carryinitout(bfn_22_21_0_));
    defparam IN_MUX_bfv_22_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_22_0_ (
            .carryinitin(un2_cntdiv_1_cry_16),
            .carryinitout(bfn_22_22_0_));
    defparam IN_MUX_bfv_22_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_23_0_ (
            .carryinitin(un2_cntdiv_1_cry_24),
            .carryinitout(bfn_22_23_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam cntDiv_1_LC_21_20_0.C_ON=1'b0;
    defparam cntDiv_1_LC_21_20_0.SEQ_MODE=4'b1000;
    defparam cntDiv_1_LC_21_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 cntDiv_1_LC_21_20_0 (
            .in0(_gnd_net_),
            .in1(N__1199),
            .in2(_gnd_net_),
            .in3(N__1175),
            .lcout(cntDivZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1580),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_0_LC_21_20_1.C_ON=1'b0;
    defparam cntDiv_0_LC_21_20_1.SEQ_MODE=4'b1000;
    defparam cntDiv_0_LC_21_20_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 cntDiv_0_LC_21_20_1 (
            .in0(N__1200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cntDivZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1580),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_cry_1_c_LC_22_17_0.C_ON=1'b1;
    defparam un2_cntdiv_cry_1_c_LC_22_17_0.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_cry_1_c_LC_22_17_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_cry_1_c_LC_22_17_0 (
            .in0(_gnd_net_),
            .in1(N__1177),
            .in2(N__1204),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_17_0_),
            .carryout(un2_cntdiv_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_2_LC_22_17_1.C_ON=1'b1;
    defparam cntDiv_2_LC_22_17_1.SEQ_MODE=4'b1000;
    defparam cntDiv_2_LC_22_17_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_2_LC_22_17_1 (
            .in0(_gnd_net_),
            .in1(N__1149),
            .in2(_gnd_net_),
            .in3(N__994),
            .lcout(cntDivZ0Z_2),
            .ltout(),
            .carryin(un2_cntdiv_cry_1),
            .carryout(un2_cntdiv_cry_2),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_3_LC_22_17_2.C_ON=1'b1;
    defparam cntDiv_3_LC_22_17_2.SEQ_MODE=4'b1000;
    defparam cntDiv_3_LC_22_17_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_3_LC_22_17_2 (
            .in0(_gnd_net_),
            .in1(N__1134),
            .in2(_gnd_net_),
            .in3(N__991),
            .lcout(cntDivZ0Z_3),
            .ltout(),
            .carryin(un2_cntdiv_cry_2),
            .carryout(un2_cntdiv_cry_3),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_4_LC_22_17_3.C_ON=1'b1;
    defparam cntDiv_4_LC_22_17_3.SEQ_MODE=4'b1000;
    defparam cntDiv_4_LC_22_17_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_4_LC_22_17_3 (
            .in0(_gnd_net_),
            .in1(N__1116),
            .in2(_gnd_net_),
            .in3(N__988),
            .lcout(cntDivZ0Z_4),
            .ltout(),
            .carryin(un2_cntdiv_cry_3),
            .carryout(un2_cntdiv_cry_4),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_5_LC_22_17_4.C_ON=1'b1;
    defparam cntDiv_5_LC_22_17_4.SEQ_MODE=4'b1000;
    defparam cntDiv_5_LC_22_17_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_5_LC_22_17_4 (
            .in0(_gnd_net_),
            .in1(N__1098),
            .in2(_gnd_net_),
            .in3(N__1021),
            .lcout(cntDivZ0Z_5),
            .ltout(),
            .carryin(un2_cntdiv_cry_4),
            .carryout(un2_cntdiv_cry_5),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_6_LC_22_17_5.C_ON=1'b1;
    defparam cntDiv_6_LC_22_17_5.SEQ_MODE=4'b1000;
    defparam cntDiv_6_LC_22_17_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_6_LC_22_17_5 (
            .in0(_gnd_net_),
            .in1(N__1080),
            .in2(_gnd_net_),
            .in3(N__1018),
            .lcout(cntDivZ0Z_6),
            .ltout(),
            .carryin(un2_cntdiv_cry_5),
            .carryout(un2_cntdiv_cry_6),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_7_LC_22_17_6.C_ON=1'b1;
    defparam cntDiv_7_LC_22_17_6.SEQ_MODE=4'b1000;
    defparam cntDiv_7_LC_22_17_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_7_LC_22_17_6 (
            .in0(_gnd_net_),
            .in1(N__1062),
            .in2(_gnd_net_),
            .in3(N__1015),
            .lcout(cntDivZ0Z_7),
            .ltout(),
            .carryin(un2_cntdiv_cry_6),
            .carryout(un2_cntdiv_cry_7),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_8_LC_22_17_7.C_ON=1'b1;
    defparam cntDiv_8_LC_22_17_7.SEQ_MODE=4'b1000;
    defparam cntDiv_8_LC_22_17_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_8_LC_22_17_7 (
            .in0(_gnd_net_),
            .in1(N__1347),
            .in2(_gnd_net_),
            .in3(N__1012),
            .lcout(cntDivZ0Z_8),
            .ltout(),
            .carryin(un2_cntdiv_cry_7),
            .carryout(un2_cntdiv_cry_8),
            .clk(N__1578),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_9_LC_22_18_0.C_ON=1'b1;
    defparam cntDiv_9_LC_22_18_0.SEQ_MODE=4'b1000;
    defparam cntDiv_9_LC_22_18_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_9_LC_22_18_0 (
            .in0(_gnd_net_),
            .in1(N__1329),
            .in2(_gnd_net_),
            .in3(N__1009),
            .lcout(cntDivZ0Z_9),
            .ltout(),
            .carryin(bfn_22_18_0_),
            .carryout(un2_cntdiv_cry_9),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_10_LC_22_18_1.C_ON=1'b1;
    defparam cntDiv_10_LC_22_18_1.SEQ_MODE=4'b1000;
    defparam cntDiv_10_LC_22_18_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_10_LC_22_18_1 (
            .in0(_gnd_net_),
            .in1(N__1311),
            .in2(_gnd_net_),
            .in3(N__1006),
            .lcout(cntDivZ0Z_10),
            .ltout(),
            .carryin(un2_cntdiv_cry_9),
            .carryout(un2_cntdiv_cry_10),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_11_LC_22_18_2.C_ON=1'b1;
    defparam cntDiv_11_LC_22_18_2.SEQ_MODE=4'b1000;
    defparam cntDiv_11_LC_22_18_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_11_LC_22_18_2 (
            .in0(_gnd_net_),
            .in1(N__1293),
            .in2(_gnd_net_),
            .in3(N__1003),
            .lcout(cntDivZ0Z_11),
            .ltout(),
            .carryin(un2_cntdiv_cry_10),
            .carryout(un2_cntdiv_cry_11),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_12_LC_22_18_3.C_ON=1'b1;
    defparam cntDiv_12_LC_22_18_3.SEQ_MODE=4'b1000;
    defparam cntDiv_12_LC_22_18_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_12_LC_22_18_3 (
            .in0(_gnd_net_),
            .in1(N__1278),
            .in2(_gnd_net_),
            .in3(N__1000),
            .lcout(cntDivZ0Z_12),
            .ltout(),
            .carryin(un2_cntdiv_cry_11),
            .carryout(un2_cntdiv_cry_12),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_13_LC_22_18_4.C_ON=1'b1;
    defparam cntDiv_13_LC_22_18_4.SEQ_MODE=4'b1000;
    defparam cntDiv_13_LC_22_18_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_13_LC_22_18_4 (
            .in0(_gnd_net_),
            .in1(N__1260),
            .in2(_gnd_net_),
            .in3(N__997),
            .lcout(cntDivZ0Z_13),
            .ltout(),
            .carryin(un2_cntdiv_cry_12),
            .carryout(un2_cntdiv_cry_13),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_14_LC_22_18_5.C_ON=1'b1;
    defparam cntDiv_14_LC_22_18_5.SEQ_MODE=4'b1000;
    defparam cntDiv_14_LC_22_18_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_14_LC_22_18_5 (
            .in0(_gnd_net_),
            .in1(N__1242),
            .in2(_gnd_net_),
            .in3(N__1048),
            .lcout(cntDivZ0Z_14),
            .ltout(),
            .carryin(un2_cntdiv_cry_13),
            .carryout(un2_cntdiv_cry_14),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_15_LC_22_18_6.C_ON=1'b1;
    defparam cntDiv_15_LC_22_18_6.SEQ_MODE=4'b1000;
    defparam cntDiv_15_LC_22_18_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_15_LC_22_18_6 (
            .in0(_gnd_net_),
            .in1(N__1224),
            .in2(_gnd_net_),
            .in3(N__1045),
            .lcout(cntDivZ0Z_15),
            .ltout(),
            .carryin(un2_cntdiv_cry_14),
            .carryout(un2_cntdiv_cry_15),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_16_LC_22_18_7.C_ON=1'b1;
    defparam cntDiv_16_LC_22_18_7.SEQ_MODE=4'b1000;
    defparam cntDiv_16_LC_22_18_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_16_LC_22_18_7 (
            .in0(_gnd_net_),
            .in1(N__1506),
            .in2(_gnd_net_),
            .in3(N__1042),
            .lcout(cntDivZ0Z_16),
            .ltout(),
            .carryin(un2_cntdiv_cry_15),
            .carryout(un2_cntdiv_cry_16),
            .clk(N__1579),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_17_LC_22_19_0.C_ON=1'b1;
    defparam cntDiv_17_LC_22_19_0.SEQ_MODE=4'b1000;
    defparam cntDiv_17_LC_22_19_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_17_LC_22_19_0 (
            .in0(_gnd_net_),
            .in1(N__1488),
            .in2(_gnd_net_),
            .in3(N__1039),
            .lcout(cntDivZ0Z_17),
            .ltout(),
            .carryin(bfn_22_19_0_),
            .carryout(un2_cntdiv_cry_17),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_18_LC_22_19_1.C_ON=1'b1;
    defparam cntDiv_18_LC_22_19_1.SEQ_MODE=4'b1000;
    defparam cntDiv_18_LC_22_19_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_18_LC_22_19_1 (
            .in0(_gnd_net_),
            .in1(N__1470),
            .in2(_gnd_net_),
            .in3(N__1036),
            .lcout(cntDivZ0Z_18),
            .ltout(),
            .carryin(un2_cntdiv_cry_17),
            .carryout(un2_cntdiv_cry_18),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_19_LC_22_19_2.C_ON=1'b1;
    defparam cntDiv_19_LC_22_19_2.SEQ_MODE=4'b1000;
    defparam cntDiv_19_LC_22_19_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_19_LC_22_19_2 (
            .in0(_gnd_net_),
            .in1(N__1452),
            .in2(_gnd_net_),
            .in3(N__1033),
            .lcout(cntDivZ0Z_19),
            .ltout(),
            .carryin(un2_cntdiv_cry_18),
            .carryout(un2_cntdiv_cry_19),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_20_LC_22_19_3.C_ON=1'b1;
    defparam cntDiv_20_LC_22_19_3.SEQ_MODE=4'b1000;
    defparam cntDiv_20_LC_22_19_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_20_LC_22_19_3 (
            .in0(_gnd_net_),
            .in1(N__1434),
            .in2(_gnd_net_),
            .in3(N__1030),
            .lcout(cntDivZ0Z_20),
            .ltout(),
            .carryin(un2_cntdiv_cry_19),
            .carryout(un2_cntdiv_cry_20),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_21_LC_22_19_4.C_ON=1'b1;
    defparam cntDiv_21_LC_22_19_4.SEQ_MODE=4'b1000;
    defparam cntDiv_21_LC_22_19_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_21_LC_22_19_4 (
            .in0(_gnd_net_),
            .in1(N__1416),
            .in2(_gnd_net_),
            .in3(N__1027),
            .lcout(cntDivZ0Z_21),
            .ltout(),
            .carryin(un2_cntdiv_cry_20),
            .carryout(un2_cntdiv_cry_21),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_22_LC_22_19_5.C_ON=1'b1;
    defparam cntDiv_22_LC_22_19_5.SEQ_MODE=4'b1000;
    defparam cntDiv_22_LC_22_19_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_22_LC_22_19_5 (
            .in0(_gnd_net_),
            .in1(N__1398),
            .in2(_gnd_net_),
            .in3(N__1024),
            .lcout(cntDivZ0Z_22),
            .ltout(),
            .carryin(un2_cntdiv_cry_21),
            .carryout(un2_cntdiv_cry_22),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_23_LC_22_19_6.C_ON=1'b1;
    defparam cntDiv_23_LC_22_19_6.SEQ_MODE=4'b1000;
    defparam cntDiv_23_LC_22_19_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntDiv_23_LC_22_19_6 (
            .in0(_gnd_net_),
            .in1(N__1380),
            .in2(_gnd_net_),
            .in3(N__1210),
            .lcout(cntDivZ0Z_23),
            .ltout(),
            .carryin(un2_cntdiv_cry_22),
            .carryout(un2_cntdiv_cry_23),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_24_LC_22_19_7.C_ON=1'b0;
    defparam cntDiv_24_LC_22_19_7.SEQ_MODE=4'b1000;
    defparam cntDiv_24_LC_22_19_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 cntDiv_24_LC_22_19_7 (
            .in0(_gnd_net_),
            .in1(N__1365),
            .in2(_gnd_net_),
            .in3(N__1207),
            .lcout(cntDivZ0Z_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1581),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_1_c_LC_22_20_0.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_1_c_LC_22_20_0.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_1_c_LC_22_20_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_1_c_LC_22_20_0 (
            .in0(_gnd_net_),
            .in1(N__1195),
            .in2(N__1176),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_20_0_),
            .carryout(un2_cntdiv_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_2_c_LC_22_20_1.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_2_c_LC_22_20_1.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_2_c_LC_22_20_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_2_c_LC_22_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1153),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_1),
            .carryout(un2_cntdiv_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_3_c_LC_22_20_2.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_3_c_LC_22_20_2.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_3_c_LC_22_20_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_3_c_LC_22_20_2 (
            .in0(_gnd_net_),
            .in1(N__1135),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_2),
            .carryout(un2_cntdiv_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_4_c_LC_22_20_3.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_4_c_LC_22_20_3.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_4_c_LC_22_20_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_4_c_LC_22_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_3),
            .carryout(un2_cntdiv_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_5_c_LC_22_20_4.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_5_c_LC_22_20_4.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_5_c_LC_22_20_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_5_c_LC_22_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1102),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_4),
            .carryout(un2_cntdiv_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_6_c_LC_22_20_5.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_6_c_LC_22_20_5.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_6_c_LC_22_20_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_6_c_LC_22_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1084),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_5),
            .carryout(un2_cntdiv_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_7_c_LC_22_20_6.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_7_c_LC_22_20_6.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_7_c_LC_22_20_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_7_c_LC_22_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1066),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_6),
            .carryout(un2_cntdiv_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_8_c_LC_22_20_7.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_8_c_LC_22_20_7.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_8_c_LC_22_20_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_8_c_LC_22_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1351),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_7),
            .carryout(un2_cntdiv_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_9_c_LC_22_21_0.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_9_c_LC_22_21_0.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_9_c_LC_22_21_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_9_c_LC_22_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1333),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_21_0_),
            .carryout(un2_cntdiv_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_10_c_LC_22_21_1.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_10_c_LC_22_21_1.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_10_c_LC_22_21_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_10_c_LC_22_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1315),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_9),
            .carryout(un2_cntdiv_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_11_c_LC_22_21_2.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_11_c_LC_22_21_2.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_11_c_LC_22_21_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_11_c_LC_22_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1297),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_10),
            .carryout(un2_cntdiv_1_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_12_c_LC_22_21_3.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_12_c_LC_22_21_3.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_12_c_LC_22_21_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_12_c_LC_22_21_3 (
            .in0(_gnd_net_),
            .in1(N__1279),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_11),
            .carryout(un2_cntdiv_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_13_c_LC_22_21_4.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_13_c_LC_22_21_4.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_13_c_LC_22_21_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_13_c_LC_22_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1264),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_12),
            .carryout(un2_cntdiv_1_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_14_c_LC_22_21_5.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_14_c_LC_22_21_5.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_14_c_LC_22_21_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_14_c_LC_22_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1246),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_13),
            .carryout(un2_cntdiv_1_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_15_c_LC_22_21_6.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_15_c_LC_22_21_6.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_15_c_LC_22_21_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_15_c_LC_22_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1228),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_14),
            .carryout(un2_cntdiv_1_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_16_c_LC_22_21_7.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_16_c_LC_22_21_7.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_16_c_LC_22_21_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_16_c_LC_22_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1510),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_15),
            .carryout(un2_cntdiv_1_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_17_c_LC_22_22_0.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_17_c_LC_22_22_0.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_17_c_LC_22_22_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_17_c_LC_22_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1492),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_22_0_),
            .carryout(un2_cntdiv_1_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_18_c_LC_22_22_1.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_18_c_LC_22_22_1.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_18_c_LC_22_22_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_18_c_LC_22_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1474),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_17),
            .carryout(un2_cntdiv_1_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_19_c_LC_22_22_2.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_19_c_LC_22_22_2.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_19_c_LC_22_22_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_19_c_LC_22_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1456),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_18),
            .carryout(un2_cntdiv_1_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_20_c_LC_22_22_3.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_20_c_LC_22_22_3.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_20_c_LC_22_22_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_20_c_LC_22_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1438),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_19),
            .carryout(un2_cntdiv_1_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_21_c_LC_22_22_4.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_21_c_LC_22_22_4.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_21_c_LC_22_22_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_21_c_LC_22_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1420),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_20),
            .carryout(un2_cntdiv_1_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_22_c_LC_22_22_5.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_22_c_LC_22_22_5.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_22_c_LC_22_22_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_22_c_LC_22_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1402),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_21),
            .carryout(un2_cntdiv_1_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_23_c_LC_22_22_6.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_23_c_LC_22_22_6.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_23_c_LC_22_22_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_23_c_LC_22_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1384),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_22),
            .carryout(un2_cntdiv_1_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_24_c_LC_22_22_7.C_ON=1'b1;
    defparam un2_cntdiv_1_cry_24_c_LC_22_22_7.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_24_c_LC_22_22_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_cntdiv_1_cry_24_c_LC_22_22_7 (
            .in0(_gnd_net_),
            .in1(N__1366),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un2_cntdiv_1_cry_23),
            .carryout(un2_cntdiv_1_cry_24),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_cntdiv_1_cry_24_c_RNI73PB_LC_22_23_0.C_ON=1'b0;
    defparam un2_cntdiv_1_cry_24_c_RNI73PB_LC_22_23_0.SEQ_MODE=4'b0000;
    defparam un2_cntdiv_1_cry_24_c_RNI73PB_LC_22_23_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 un2_cntdiv_1_cry_24_c_RNI73PB_LC_22_23_0 (
            .in0(_gnd_net_),
            .in1(N__1596),
            .in2(_gnd_net_),
            .in3(N__1612),
            .lcout(un2_cntdiv_1_cry_24_c_RNI73PBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \counter1.Pre_Q_1_LC_23_21_5 .C_ON=1'b0;
    defparam \counter1.Pre_Q_1_LC_23_21_5 .SEQ_MODE=4'b1000;
    defparam \counter1.Pre_Q_1_LC_23_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \counter1.Pre_Q_1_LC_23_21_5  (
            .in0(N__1811),
            .in1(N__1879),
            .in2(_gnd_net_),
            .in3(N__1678),
            .lcout(value_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1582),
            .ce(N__1551),
            .sr(_gnd_net_));
    defparam cntDiv_RNIETOH_25_LC_23_22_4.C_ON=1'b0;
    defparam cntDiv_RNIETOH_25_LC_23_22_4.SEQ_MODE=4'b0000;
    defparam cntDiv_RNIETOH_25_LC_23_22_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 cntDiv_RNIETOH_25_LC_23_22_4 (
            .in0(_gnd_net_),
            .in1(N__1597),
            .in2(_gnd_net_),
            .in3(N__1608),
            .lcout(cntDiv_RNIETOHZ0Z_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntDiv_25_LC_23_23_1.C_ON=1'b0;
    defparam cntDiv_25_LC_23_23_1.SEQ_MODE=4'b1000;
    defparam cntDiv_25_LC_23_23_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 cntDiv_25_LC_23_23_1 (
            .in0(_gnd_net_),
            .in1(N__1609),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cntDiv_i_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1584),
            .ce(),
            .sr(_gnd_net_));
    defparam \counter1.Pre_Q_3_LC_24_21_4 .C_ON=1'b0;
    defparam \counter1.Pre_Q_3_LC_24_21_4 .SEQ_MODE=4'b1000;
    defparam \counter1.Pre_Q_3_LC_24_21_4 .LUT_INIT=16'b0100000000000010;
    LogicCell40 \counter1.Pre_Q_3_LC_24_21_4  (
            .in0(N__1812),
            .in1(N__1880),
            .in2(N__1691),
            .in3(N__1741),
            .lcout(value_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1583),
            .ce(N__1555),
            .sr(_gnd_net_));
    defparam \counter1.Pre_Q_2_LC_24_22_2 .C_ON=1'b0;
    defparam \counter1.Pre_Q_2_LC_24_22_2 .SEQ_MODE=4'b1000;
    defparam \counter1.Pre_Q_2_LC_24_22_2 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \counter1.Pre_Q_2_LC_24_22_2  (
            .in0(N__1673),
            .in1(N__1814),
            .in2(N__1898),
            .in3(N__1740),
            .lcout(value_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1585),
            .ce(N__1550),
            .sr(_gnd_net_));
    defparam \counter1.Pre_Q_0_LC_24_22_7 .C_ON=1'b0;
    defparam \counter1.Pre_Q_0_LC_24_22_7 .SEQ_MODE=4'b1000;
    defparam \counter1.Pre_Q_0_LC_24_22_7 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \counter1.Pre_Q_0_LC_24_22_7  (
            .in0(N__1813),
            .in1(N__1881),
            .in2(N__1748),
            .in3(N__1674),
            .lcout(value_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__1585),
            .ce(N__1550),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m6_LC_32_21_0 .C_ON=1'b0;
    defparam \display.S_1_7_0__m6_LC_32_21_0 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m6_LC_32_21_0 .LUT_INIT=16'b0001001101100110;
    LogicCell40 \display.S_1_7_0__m6_LC_32_21_0  (
            .in0(N__1783),
            .in1(N__1830),
            .in2(N__1714),
            .in3(N__1903),
            .lcout(Y_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m15_LC_32_21_4 .C_ON=1'b0;
    defparam \display.S_1_7_0__m15_LC_32_21_4 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m15_LC_32_21_4 .LUT_INIT=16'b0001001100100100;
    LogicCell40 \display.S_1_7_0__m15_LC_32_21_4  (
            .in0(N__1781),
            .in1(N__1828),
            .in2(N__1713),
            .in3(N__1902),
            .lcout(Y_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m2_LC_32_21_5 .C_ON=1'b0;
    defparam \display.S_1_7_0__m2_LC_32_21_5 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m2_LC_32_21_5 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \display.S_1_7_0__m2_LC_32_21_5  (
            .in0(N__1829),
            .in1(N__1782),
            .in2(_gnd_net_),
            .in3(N__1904),
            .lcout(Y_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m11_LC_32_21_7 .C_ON=1'b0;
    defparam \display.S_1_7_0__m11_LC_32_21_7 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m11_LC_32_21_7 .LUT_INIT=16'b0000011001000110;
    LogicCell40 \display.S_1_7_0__m11_LC_32_21_7  (
            .in0(N__1827),
            .in1(N__1780),
            .in2(N__1908),
            .in3(N__1706),
            .lcout(Y_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m19_LC_32_22_0 .C_ON=1'b0;
    defparam \display.S_1_7_0__m19_LC_32_22_0 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m19_LC_32_22_0 .LUT_INIT=16'b0000111100111000;
    LogicCell40 \display.S_1_7_0__m19_LC_32_22_0  (
            .in0(N__1695),
            .in1(N__1768),
            .in2(N__1852),
            .in3(N__1921),
            .lcout(Y_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m18_LC_32_22_3 .C_ON=1'b0;
    defparam \display.S_1_7_0__m18_LC_32_22_3 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m18_LC_32_22_3 .LUT_INIT=16'b0010011100010110;
    LogicCell40 \display.S_1_7_0__m18_LC_32_22_3  (
            .in0(N__1920),
            .in1(N__1847),
            .in2(N__1779),
            .in3(N__1694),
            .lcout(Y_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m13_LC_32_22_4 .C_ON=1'b0;
    defparam \display.S_1_7_0__m13_LC_32_22_4 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m13_LC_32_22_4 .LUT_INIT=16'b0000010100010000;
    LogicCell40 \display.S_1_7_0__m13_LC_32_22_4  (
            .in0(N__1692),
            .in1(N__1761),
            .in2(N__1851),
            .in3(N__1918),
            .lcout(Y_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \display.S_1_7_0__m16_LC_32_22_5 .C_ON=1'b0;
    defparam \display.S_1_7_0__m16_LC_32_22_5 .SEQ_MODE=4'b0000;
    defparam \display.S_1_7_0__m16_LC_32_22_5 .LUT_INIT=16'b0011011100110100;
    LogicCell40 \display.S_1_7_0__m16_LC_32_22_5  (
            .in0(N__1919),
            .in1(N__1846),
            .in2(N__1778),
            .in3(N__1693),
            .lcout(Y_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_32_28_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_32_28_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_32_28_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_32_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
