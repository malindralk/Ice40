-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 15 2022 06:07:59

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    Y : out std_logic_vector(7 downto 0);
    mclock : in std_logic;
    DIGIT1 : out std_logic;
    DIGIT2 : out std_logic;
    DIGIT3 : out std_logic;
    DIGIT4 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__2101\ : std_logic;
signal \N__2100\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2088\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2052\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2036\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2025\ : std_logic;
signal \N__2018\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2008\ : std_logic;
signal \N__2007\ : std_logic;
signal \N__2000\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1972\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1948\ : std_logic;
signal \N__1945\ : std_logic;
signal \N__1942\ : std_logic;
signal \N__1939\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1924\ : std_logic;
signal \N__1921\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1909\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1902\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1848\ : std_logic;
signal \N__1847\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1834\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1830\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1827\ : std_logic;
signal \N__1824\ : std_logic;
signal \N__1815\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1812\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1800\ : std_logic;
signal \N__1797\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1782\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1779\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1749\ : std_logic;
signal \N__1748\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1742\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1734\ : std_logic;
signal \N__1731\ : std_logic;
signal \N__1728\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1694\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1691\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1679\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1674\ : std_logic;
signal \N__1673\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1636\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1624\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1608\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1590\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1583\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1581\ : std_logic;
signal \N__1580\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1578\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1558\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1551\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1547\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1500\ : std_logic;
signal \N__1497\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1488\ : std_logic;
signal \N__1485\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1479\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1467\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1452\ : std_logic;
signal \N__1449\ : std_logic;
signal \N__1446\ : std_logic;
signal \N__1443\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1435\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1431\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1420\ : std_logic;
signal \N__1417\ : std_logic;
signal \N__1416\ : std_logic;
signal \N__1413\ : std_logic;
signal \N__1410\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1398\ : std_logic;
signal \N__1395\ : std_logic;
signal \N__1392\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1384\ : std_logic;
signal \N__1381\ : std_logic;
signal \N__1380\ : std_logic;
signal \N__1377\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1366\ : std_logic;
signal \N__1365\ : std_logic;
signal \N__1362\ : std_logic;
signal \N__1359\ : std_logic;
signal \N__1356\ : std_logic;
signal \N__1351\ : std_logic;
signal \N__1348\ : std_logic;
signal \N__1347\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1341\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1333\ : std_logic;
signal \N__1330\ : std_logic;
signal \N__1329\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1323\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1315\ : std_logic;
signal \N__1312\ : std_logic;
signal \N__1311\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1302\ : std_logic;
signal \N__1297\ : std_logic;
signal \N__1294\ : std_logic;
signal \N__1293\ : std_logic;
signal \N__1290\ : std_logic;
signal \N__1287\ : std_logic;
signal \N__1284\ : std_logic;
signal \N__1279\ : std_logic;
signal \N__1278\ : std_logic;
signal \N__1275\ : std_logic;
signal \N__1272\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1264\ : std_logic;
signal \N__1261\ : std_logic;
signal \N__1260\ : std_logic;
signal \N__1257\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1246\ : std_logic;
signal \N__1243\ : std_logic;
signal \N__1242\ : std_logic;
signal \N__1239\ : std_logic;
signal \N__1236\ : std_logic;
signal \N__1233\ : std_logic;
signal \N__1228\ : std_logic;
signal \N__1225\ : std_logic;
signal \N__1224\ : std_logic;
signal \N__1221\ : std_logic;
signal \N__1218\ : std_logic;
signal \N__1215\ : std_logic;
signal \N__1210\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1204\ : std_logic;
signal \N__1201\ : std_logic;
signal \N__1200\ : std_logic;
signal \N__1199\ : std_logic;
signal \N__1196\ : std_logic;
signal \N__1195\ : std_logic;
signal \N__1190\ : std_logic;
signal \N__1187\ : std_logic;
signal \N__1184\ : std_logic;
signal \N__1177\ : std_logic;
signal \N__1176\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1172\ : std_logic;
signal \N__1169\ : std_logic;
signal \N__1166\ : std_logic;
signal \N__1163\ : std_logic;
signal \N__1160\ : std_logic;
signal \N__1153\ : std_logic;
signal \N__1150\ : std_logic;
signal \N__1149\ : std_logic;
signal \N__1146\ : std_logic;
signal \N__1143\ : std_logic;
signal \N__1140\ : std_logic;
signal \N__1135\ : std_logic;
signal \N__1134\ : std_logic;
signal \N__1131\ : std_logic;
signal \N__1128\ : std_logic;
signal \N__1125\ : std_logic;
signal \N__1120\ : std_logic;
signal \N__1117\ : std_logic;
signal \N__1116\ : std_logic;
signal \N__1113\ : std_logic;
signal \N__1110\ : std_logic;
signal \N__1107\ : std_logic;
signal \N__1102\ : std_logic;
signal \N__1099\ : std_logic;
signal \N__1098\ : std_logic;
signal \N__1095\ : std_logic;
signal \N__1092\ : std_logic;
signal \N__1089\ : std_logic;
signal \N__1084\ : std_logic;
signal \N__1081\ : std_logic;
signal \N__1080\ : std_logic;
signal \N__1077\ : std_logic;
signal \N__1074\ : std_logic;
signal \N__1071\ : std_logic;
signal \N__1066\ : std_logic;
signal \N__1063\ : std_logic;
signal \N__1062\ : std_logic;
signal \N__1059\ : std_logic;
signal \N__1056\ : std_logic;
signal \N__1053\ : std_logic;
signal \N__1048\ : std_logic;
signal \N__1045\ : std_logic;
signal \N__1042\ : std_logic;
signal \N__1039\ : std_logic;
signal \N__1036\ : std_logic;
signal \N__1033\ : std_logic;
signal \N__1030\ : std_logic;
signal \N__1027\ : std_logic;
signal \N__1024\ : std_logic;
signal \N__1021\ : std_logic;
signal \N__1018\ : std_logic;
signal \N__1015\ : std_logic;
signal \N__1012\ : std_logic;
signal \N__1009\ : std_logic;
signal \N__1006\ : std_logic;
signal \N__1003\ : std_logic;
signal \N__1000\ : std_logic;
signal \N__997\ : std_logic;
signal \N__994\ : std_logic;
signal \N__991\ : std_logic;
signal \N__988\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_22_17_0_\ : std_logic;
signal un2_cntdiv_cry_1 : std_logic;
signal un2_cntdiv_cry_2 : std_logic;
signal un2_cntdiv_cry_3 : std_logic;
signal un2_cntdiv_cry_4 : std_logic;
signal un2_cntdiv_cry_5 : std_logic;
signal un2_cntdiv_cry_6 : std_logic;
signal un2_cntdiv_cry_7 : std_logic;
signal un2_cntdiv_cry_8 : std_logic;
signal \bfn_22_18_0_\ : std_logic;
signal un2_cntdiv_cry_9 : std_logic;
signal un2_cntdiv_cry_10 : std_logic;
signal un2_cntdiv_cry_11 : std_logic;
signal un2_cntdiv_cry_12 : std_logic;
signal un2_cntdiv_cry_13 : std_logic;
signal un2_cntdiv_cry_14 : std_logic;
signal un2_cntdiv_cry_15 : std_logic;
signal un2_cntdiv_cry_16 : std_logic;
signal \bfn_22_19_0_\ : std_logic;
signal un2_cntdiv_cry_17 : std_logic;
signal un2_cntdiv_cry_18 : std_logic;
signal un2_cntdiv_cry_19 : std_logic;
signal un2_cntdiv_cry_20 : std_logic;
signal un2_cntdiv_cry_21 : std_logic;
signal un2_cntdiv_cry_22 : std_logic;
signal un2_cntdiv_cry_23 : std_logic;
signal \cntDivZ0Z_0\ : std_logic;
signal \cntDivZ0Z_1\ : std_logic;
signal \bfn_22_20_0_\ : std_logic;
signal \cntDivZ0Z_2\ : std_logic;
signal un2_cntdiv_1_cry_1 : std_logic;
signal \cntDivZ0Z_3\ : std_logic;
signal un2_cntdiv_1_cry_2 : std_logic;
signal \cntDivZ0Z_4\ : std_logic;
signal un2_cntdiv_1_cry_3 : std_logic;
signal \cntDivZ0Z_5\ : std_logic;
signal un2_cntdiv_1_cry_4 : std_logic;
signal \cntDivZ0Z_6\ : std_logic;
signal un2_cntdiv_1_cry_5 : std_logic;
signal \cntDivZ0Z_7\ : std_logic;
signal un2_cntdiv_1_cry_6 : std_logic;
signal \cntDivZ0Z_8\ : std_logic;
signal un2_cntdiv_1_cry_7 : std_logic;
signal un2_cntdiv_1_cry_8 : std_logic;
signal \cntDivZ0Z_9\ : std_logic;
signal \bfn_22_21_0_\ : std_logic;
signal \cntDivZ0Z_10\ : std_logic;
signal un2_cntdiv_1_cry_9 : std_logic;
signal \cntDivZ0Z_11\ : std_logic;
signal un2_cntdiv_1_cry_10 : std_logic;
signal \cntDivZ0Z_12\ : std_logic;
signal un2_cntdiv_1_cry_11 : std_logic;
signal \cntDivZ0Z_13\ : std_logic;
signal un2_cntdiv_1_cry_12 : std_logic;
signal \cntDivZ0Z_14\ : std_logic;
signal un2_cntdiv_1_cry_13 : std_logic;
signal \cntDivZ0Z_15\ : std_logic;
signal un2_cntdiv_1_cry_14 : std_logic;
signal \cntDivZ0Z_16\ : std_logic;
signal un2_cntdiv_1_cry_15 : std_logic;
signal un2_cntdiv_1_cry_16 : std_logic;
signal \cntDivZ0Z_17\ : std_logic;
signal \bfn_22_22_0_\ : std_logic;
signal \cntDivZ0Z_18\ : std_logic;
signal un2_cntdiv_1_cry_17 : std_logic;
signal \cntDivZ0Z_19\ : std_logic;
signal un2_cntdiv_1_cry_18 : std_logic;
signal \cntDivZ0Z_20\ : std_logic;
signal un2_cntdiv_1_cry_19 : std_logic;
signal \cntDivZ0Z_21\ : std_logic;
signal un2_cntdiv_1_cry_20 : std_logic;
signal \cntDivZ0Z_22\ : std_logic;
signal un2_cntdiv_1_cry_21 : std_logic;
signal \cntDivZ0Z_23\ : std_logic;
signal un2_cntdiv_1_cry_22 : std_logic;
signal \cntDivZ0Z_24\ : std_logic;
signal un2_cntdiv_1_cry_23 : std_logic;
signal un2_cntdiv_1_cry_24 : std_logic;
signal \bfn_22_23_0_\ : std_logic;
signal \un2_cntdiv_1_cry_24_c_RNI73PBZ0\ : std_logic;
signal \cntDiv_i_25\ : std_logic;
signal mclock_0_c_g : std_logic;
signal \cntDiv_RNIETOHZ0Z_25\ : std_logic;
signal \Y_c_1\ : std_logic;
signal \Y_c_4\ : std_logic;
signal \Y_c_0\ : std_logic;
signal \Y_c_2\ : std_logic;
signal \Y_c_7\ : std_logic;
signal \Y_c_6\ : std_logic;
signal \Y_c_3\ : std_logic;
signal value_1 : std_logic;
signal value_3 : std_logic;
signal value_2 : std_logic;
signal value_0 : std_logic;
signal \Y_c_5\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal mclock_wire : std_logic;
signal \Y_wire\ : std_logic_vector(7 downto 0);
signal \DIGIT2_wire\ : std_logic;
signal \DIGIT1_wire\ : std_logic;
signal \DIGIT3_wire\ : std_logic;
signal \DIGIT4_wire\ : std_logic;

begin
    mclock_wire <= mclock;
    Y <= \Y_wire\;
    DIGIT2 <= \DIGIT2_wire\;
    DIGIT1 <= \DIGIT1_wire\;
    DIGIT3 <= \DIGIT3_wire\;
    DIGIT4 <= \DIGIT4_wire\;

    \mclock_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2099\,
            GLOBALBUFFEROUTPUT => mclock_0_c_g
        );

    \mclock_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2101\,
            DIN => \N__2100\,
            DOUT => \N__2099\,
            PACKAGEPIN => mclock_wire
        );

    \mclock_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2101\,
            PADOUT => \N__2100\,
            PADIN => \N__2099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2090\,
            DIN => \N__2089\,
            DOUT => \N__2088\,
            PACKAGEPIN => \Y_wire\(7)
        );

    \Y_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2090\,
            PADOUT => \N__2089\,
            PADIN => \N__2088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1948\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2081\,
            DIN => \N__2080\,
            DOUT => \N__2079\,
            PACKAGEPIN => \Y_wire\(0)
        );

    \Y_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2081\,
            PADOUT => \N__2080\,
            PADIN => \N__2079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1972\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DIGIT2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2072\,
            DIN => \N__2071\,
            DOUT => \N__2070\,
            PACKAGEPIN => \DIGIT2_wire\
        );

    \DIGIT2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2072\,
            PADOUT => \N__2071\,
            PADIN => \N__2070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2063\,
            DIN => \N__2062\,
            DOUT => \N__2061\,
            PACKAGEPIN => \Y_wire\(4)
        );

    \Y_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2063\,
            PADOUT => \N__2062\,
            PADIN => \N__2061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1516\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DIGIT1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2054\,
            DIN => \N__2053\,
            DOUT => \N__2052\,
            PACKAGEPIN => \DIGIT1_wire\
        );

    \DIGIT1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2054\,
            PADOUT => \N__2053\,
            PADIN => \N__2052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2045\,
            DIN => \N__2044\,
            DOUT => \N__2043\,
            PACKAGEPIN => \Y_wire\(1)
        );

    \Y_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2045\,
            PADOUT => \N__2044\,
            PADIN => \N__2043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1522\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2036\,
            DIN => \N__2035\,
            DOUT => \N__2034\,
            PACKAGEPIN => \Y_wire\(5)
        );

    \Y_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2036\,
            PADOUT => \N__2035\,
            PADIN => \N__2034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1645\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DIGIT3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2027\,
            DIN => \N__2026\,
            DOUT => \N__2025\,
            PACKAGEPIN => \DIGIT3_wire\
        );

    \DIGIT3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2027\,
            PADOUT => \N__2026\,
            PADIN => \N__2025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1623\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2018\,
            DIN => \N__2017\,
            DOUT => \N__2016\,
            PACKAGEPIN => \Y_wire\(2)
        );

    \Y_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2018\,
            PADOUT => \N__2017\,
            PADIN => \N__2016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1960\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DIGIT4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2009\,
            DIN => \N__2008\,
            DOUT => \N__2007\,
            PACKAGEPIN => \DIGIT4_wire\
        );

    \DIGIT4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2009\,
            PADOUT => \N__2008\,
            PADIN => \N__2007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2000\,
            DIN => \N__1999\,
            DOUT => \N__1998\,
            PACKAGEPIN => \Y_wire\(6)
        );

    \Y_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2000\,
            PADOUT => \N__1999\,
            PADIN => \N__1998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Y_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__1991\,
            DIN => \N__1990\,
            DOUT => \N__1989\,
            PACKAGEPIN => \Y_wire\(3)
        );

    \Y_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__1991\,
            PADOUT => \N__1990\,
            PADIN => \N__1989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__417\ : IoInMux
    port map (
            O => \N__1972\,
            I => \N__1969\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__1969\,
            I => \N__1966\
        );

    \I__415\ : Span4Mux_s0_h
    port map (
            O => \N__1966\,
            I => \N__1963\
        );

    \I__414\ : Odrv4
    port map (
            O => \N__1963\,
            I => \Y_c_0\
        );

    \I__413\ : IoInMux
    port map (
            O => \N__1960\,
            I => \N__1957\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__1957\,
            I => \N__1954\
        );

    \I__411\ : Span4Mux_s0_h
    port map (
            O => \N__1954\,
            I => \N__1951\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__1951\,
            I => \Y_c_2\
        );

    \I__409\ : IoInMux
    port map (
            O => \N__1948\,
            I => \N__1945\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__1945\,
            I => \N__1942\
        );

    \I__407\ : Span4Mux_s1_h
    port map (
            O => \N__1942\,
            I => \N__1939\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__1939\,
            I => \N__1936\
        );

    \I__405\ : Odrv4
    port map (
            O => \N__1936\,
            I => \Y_c_7\
        );

    \I__404\ : IoInMux
    port map (
            O => \N__1933\,
            I => \N__1930\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__1930\,
            I => \Y_c_6\
        );

    \I__402\ : IoInMux
    port map (
            O => \N__1927\,
            I => \N__1924\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__1924\,
            I => \Y_c_3\
        );

    \I__400\ : InMux
    port map (
            O => \N__1921\,
            I => \N__1909\
        );

    \I__399\ : InMux
    port map (
            O => \N__1920\,
            I => \N__1909\
        );

    \I__398\ : InMux
    port map (
            O => \N__1919\,
            I => \N__1909\
        );

    \I__397\ : InMux
    port map (
            O => \N__1918\,
            I => \N__1909\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__1909\,
            I => \N__1905\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__1908\,
            I => \N__1899\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__1905\,
            I => \N__1895\
        );

    \I__393\ : InMux
    port map (
            O => \N__1904\,
            I => \N__1892\
        );

    \I__392\ : InMux
    port map (
            O => \N__1903\,
            I => \N__1885\
        );

    \I__391\ : InMux
    port map (
            O => \N__1902\,
            I => \N__1885\
        );

    \I__390\ : InMux
    port map (
            O => \N__1899\,
            I => \N__1885\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__1898\,
            I => \N__1882\
        );

    \I__388\ : Sp12to4
    port map (
            O => \N__1895\,
            I => \N__1872\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__1892\,
            I => \N__1872\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__1885\,
            I => \N__1872\
        );

    \I__385\ : InMux
    port map (
            O => \N__1882\,
            I => \N__1867\
        );

    \I__384\ : InMux
    port map (
            O => \N__1881\,
            I => \N__1867\
        );

    \I__383\ : InMux
    port map (
            O => \N__1880\,
            I => \N__1864\
        );

    \I__382\ : InMux
    port map (
            O => \N__1879\,
            I => \N__1861\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__1872\,
            I => value_1
        );

    \I__380\ : LocalMux
    port map (
            O => \N__1867\,
            I => value_1
        );

    \I__379\ : LocalMux
    port map (
            O => \N__1864\,
            I => value_1
        );

    \I__378\ : LocalMux
    port map (
            O => \N__1861\,
            I => value_1
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__1852\,
            I => \N__1848\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__1851\,
            I => \N__1843\
        );

    \I__375\ : InMux
    port map (
            O => \N__1848\,
            I => \N__1834\
        );

    \I__374\ : InMux
    port map (
            O => \N__1847\,
            I => \N__1834\
        );

    \I__373\ : InMux
    port map (
            O => \N__1846\,
            I => \N__1834\
        );

    \I__372\ : InMux
    port map (
            O => \N__1843\,
            I => \N__1834\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__1834\,
            I => \N__1831\
        );

    \I__370\ : Span4Mux_v
    port map (
            O => \N__1831\,
            I => \N__1824\
        );

    \I__369\ : InMux
    port map (
            O => \N__1830\,
            I => \N__1815\
        );

    \I__368\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1815\
        );

    \I__367\ : InMux
    port map (
            O => \N__1828\,
            I => \N__1815\
        );

    \I__366\ : InMux
    port map (
            O => \N__1827\,
            I => \N__1815\
        );

    \I__365\ : Span4Mux_h
    port map (
            O => \N__1824\,
            I => \N__1808\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__1815\,
            I => \N__1805\
        );

    \I__363\ : InMux
    port map (
            O => \N__1814\,
            I => \N__1800\
        );

    \I__362\ : InMux
    port map (
            O => \N__1813\,
            I => \N__1800\
        );

    \I__361\ : InMux
    port map (
            O => \N__1812\,
            I => \N__1797\
        );

    \I__360\ : InMux
    port map (
            O => \N__1811\,
            I => \N__1794\
        );

    \I__359\ : Odrv4
    port map (
            O => \N__1808\,
            I => value_3
        );

    \I__358\ : Odrv12
    port map (
            O => \N__1805\,
            I => value_3
        );

    \I__357\ : LocalMux
    port map (
            O => \N__1800\,
            I => value_3
        );

    \I__356\ : LocalMux
    port map (
            O => \N__1797\,
            I => value_3
        );

    \I__355\ : LocalMux
    port map (
            O => \N__1794\,
            I => value_3
        );

    \I__354\ : InMux
    port map (
            O => \N__1783\,
            I => \N__1769\
        );

    \I__353\ : InMux
    port map (
            O => \N__1782\,
            I => \N__1769\
        );

    \I__352\ : InMux
    port map (
            O => \N__1781\,
            I => \N__1769\
        );

    \I__351\ : InMux
    port map (
            O => \N__1780\,
            I => \N__1769\
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__1779\,
            I => \N__1765\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__1778\,
            I => \N__1762\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__1769\,
            I => \N__1758\
        );

    \I__347\ : InMux
    port map (
            O => \N__1768\,
            I => \N__1749\
        );

    \I__346\ : InMux
    port map (
            O => \N__1765\,
            I => \N__1749\
        );

    \I__345\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1749\
        );

    \I__344\ : InMux
    port map (
            O => \N__1761\,
            I => \N__1749\
        );

    \I__343\ : Span4Mux_v
    port map (
            O => \N__1758\,
            I => \N__1745\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__1749\,
            I => \N__1742\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__1748\,
            I => \N__1737\
        );

    \I__340\ : Span4Mux_h
    port map (
            O => \N__1745\,
            I => \N__1734\
        );

    \I__339\ : Span12Mux_s2_h
    port map (
            O => \N__1742\,
            I => \N__1731\
        );

    \I__338\ : InMux
    port map (
            O => \N__1741\,
            I => \N__1728\
        );

    \I__337\ : InMux
    port map (
            O => \N__1740\,
            I => \N__1723\
        );

    \I__336\ : InMux
    port map (
            O => \N__1737\,
            I => \N__1723\
        );

    \I__335\ : Odrv4
    port map (
            O => \N__1734\,
            I => value_2
        );

    \I__334\ : Odrv12
    port map (
            O => \N__1731\,
            I => value_2
        );

    \I__333\ : LocalMux
    port map (
            O => \N__1728\,
            I => value_2
        );

    \I__332\ : LocalMux
    port map (
            O => \N__1723\,
            I => value_2
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__1714\,
            I => \N__1710\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__1713\,
            I => \N__1707\
        );

    \I__329\ : InMux
    port map (
            O => \N__1710\,
            I => \N__1699\
        );

    \I__328\ : InMux
    port map (
            O => \N__1707\,
            I => \N__1699\
        );

    \I__327\ : InMux
    port map (
            O => \N__1706\,
            I => \N__1699\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1699\,
            I => \N__1696\
        );

    \I__325\ : Span4Mux_s3_h
    port map (
            O => \N__1696\,
            I => \N__1688\
        );

    \I__324\ : InMux
    port map (
            O => \N__1695\,
            I => \N__1679\
        );

    \I__323\ : InMux
    port map (
            O => \N__1694\,
            I => \N__1679\
        );

    \I__322\ : InMux
    port map (
            O => \N__1693\,
            I => \N__1679\
        );

    \I__321\ : InMux
    port map (
            O => \N__1692\,
            I => \N__1679\
        );

    \I__320\ : CascadeMux
    port map (
            O => \N__1691\,
            I => \N__1675\
        );

    \I__319\ : Span4Mux_h
    port map (
            O => \N__1688\,
            I => \N__1670\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1679\,
            I => \N__1667\
        );

    \I__317\ : InMux
    port map (
            O => \N__1678\,
            I => \N__1664\
        );

    \I__316\ : InMux
    port map (
            O => \N__1675\,
            I => \N__1661\
        );

    \I__315\ : InMux
    port map (
            O => \N__1674\,
            I => \N__1656\
        );

    \I__314\ : InMux
    port map (
            O => \N__1673\,
            I => \N__1656\
        );

    \I__313\ : Odrv4
    port map (
            O => \N__1670\,
            I => value_0
        );

    \I__312\ : Odrv12
    port map (
            O => \N__1667\,
            I => value_0
        );

    \I__311\ : LocalMux
    port map (
            O => \N__1664\,
            I => value_0
        );

    \I__310\ : LocalMux
    port map (
            O => \N__1661\,
            I => value_0
        );

    \I__309\ : LocalMux
    port map (
            O => \N__1656\,
            I => value_0
        );

    \I__308\ : IoInMux
    port map (
            O => \N__1645\,
            I => \N__1642\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1642\,
            I => \N__1639\
        );

    \I__306\ : Span12Mux_s0_h
    port map (
            O => \N__1639\,
            I => \N__1636\
        );

    \I__305\ : Odrv12
    port map (
            O => \N__1636\,
            I => \Y_c_5\
        );

    \I__304\ : IoInMux
    port map (
            O => \N__1633\,
            I => \N__1630\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__1630\,
            I => \N__1627\
        );

    \I__302\ : IoSpan4Mux
    port map (
            O => \N__1627\,
            I => \N__1624\
        );

    \I__301\ : Span4Mux_s2_v
    port map (
            O => \N__1624\,
            I => \N__1620\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__1623\,
            I => \N__1617\
        );

    \I__299\ : Odrv4
    port map (
            O => \N__1620\,
            I => \CONSTANT_ONE_NET\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1617\,
            I => \CONSTANT_ONE_NET\
        );

    \I__297\ : InMux
    port map (
            O => \N__1612\,
            I => \bfn_22_23_0_\
        );

    \I__296\ : InMux
    port map (
            O => \N__1609\,
            I => \N__1605\
        );

    \I__295\ : InMux
    port map (
            O => \N__1608\,
            I => \N__1602\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1605\,
            I => \un2_cntdiv_1_cry_24_c_RNI73PBZ0\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1602\,
            I => \un2_cntdiv_1_cry_24_c_RNI73PBZ0\
        );

    \I__292\ : InMux
    port map (
            O => \N__1597\,
            I => \N__1593\
        );

    \I__291\ : InMux
    port map (
            O => \N__1596\,
            I => \N__1590\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__1593\,
            I => \cntDiv_i_25\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__1590\,
            I => \cntDiv_i_25\
        );

    \I__288\ : ClkMux
    port map (
            O => \N__1585\,
            I => \N__1561\
        );

    \I__287\ : ClkMux
    port map (
            O => \N__1584\,
            I => \N__1561\
        );

    \I__286\ : ClkMux
    port map (
            O => \N__1583\,
            I => \N__1561\
        );

    \I__285\ : ClkMux
    port map (
            O => \N__1582\,
            I => \N__1561\
        );

    \I__284\ : ClkMux
    port map (
            O => \N__1581\,
            I => \N__1561\
        );

    \I__283\ : ClkMux
    port map (
            O => \N__1580\,
            I => \N__1561\
        );

    \I__282\ : ClkMux
    port map (
            O => \N__1579\,
            I => \N__1561\
        );

    \I__281\ : ClkMux
    port map (
            O => \N__1578\,
            I => \N__1561\
        );

    \I__280\ : GlobalMux
    port map (
            O => \N__1561\,
            I => \N__1558\
        );

    \I__279\ : gio2CtrlBuf
    port map (
            O => \N__1558\,
            I => mclock_0_c_g
        );

    \I__278\ : CEMux
    port map (
            O => \N__1555\,
            I => \N__1552\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1552\,
            I => \N__1547\
        );

    \I__276\ : CEMux
    port map (
            O => \N__1551\,
            I => \N__1544\
        );

    \I__275\ : CEMux
    port map (
            O => \N__1550\,
            I => \N__1541\
        );

    \I__274\ : Span4Mux_h
    port map (
            O => \N__1547\,
            I => \N__1538\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1544\,
            I => \N__1535\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__1541\,
            I => \N__1532\
        );

    \I__271\ : Span4Mux_h
    port map (
            O => \N__1538\,
            I => \N__1527\
        );

    \I__270\ : Span4Mux_h
    port map (
            O => \N__1535\,
            I => \N__1527\
        );

    \I__269\ : Odrv12
    port map (
            O => \N__1532\,
            I => \cntDiv_RNIETOHZ0Z_25\
        );

    \I__268\ : Odrv4
    port map (
            O => \N__1527\,
            I => \cntDiv_RNIETOHZ0Z_25\
        );

    \I__267\ : IoInMux
    port map (
            O => \N__1522\,
            I => \N__1519\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1519\,
            I => \Y_c_1\
        );

    \I__265\ : IoInMux
    port map (
            O => \N__1516\,
            I => \N__1513\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1513\,
            I => \Y_c_4\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__1510\,
            I => \N__1507\
        );

    \I__262\ : InMux
    port map (
            O => \N__1507\,
            I => \N__1503\
        );

    \I__261\ : InMux
    port map (
            O => \N__1506\,
            I => \N__1500\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__1503\,
            I => \N__1497\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1500\,
            I => \cntDivZ0Z_16\
        );

    \I__258\ : Odrv4
    port map (
            O => \N__1497\,
            I => \cntDivZ0Z_16\
        );

    \I__257\ : CascadeMux
    port map (
            O => \N__1492\,
            I => \N__1489\
        );

    \I__256\ : InMux
    port map (
            O => \N__1489\,
            I => \N__1485\
        );

    \I__255\ : InMux
    port map (
            O => \N__1488\,
            I => \N__1482\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1485\,
            I => \N__1479\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__1482\,
            I => \cntDivZ0Z_17\
        );

    \I__252\ : Odrv12
    port map (
            O => \N__1479\,
            I => \cntDivZ0Z_17\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__1474\,
            I => \N__1471\
        );

    \I__250\ : InMux
    port map (
            O => \N__1471\,
            I => \N__1467\
        );

    \I__249\ : InMux
    port map (
            O => \N__1470\,
            I => \N__1464\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1467\,
            I => \N__1461\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1464\,
            I => \cntDivZ0Z_18\
        );

    \I__246\ : Odrv12
    port map (
            O => \N__1461\,
            I => \cntDivZ0Z_18\
        );

    \I__245\ : CascadeMux
    port map (
            O => \N__1456\,
            I => \N__1453\
        );

    \I__244\ : InMux
    port map (
            O => \N__1453\,
            I => \N__1449\
        );

    \I__243\ : InMux
    port map (
            O => \N__1452\,
            I => \N__1446\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1449\,
            I => \N__1443\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1446\,
            I => \cntDivZ0Z_19\
        );

    \I__240\ : Odrv4
    port map (
            O => \N__1443\,
            I => \cntDivZ0Z_19\
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__1438\,
            I => \N__1435\
        );

    \I__238\ : InMux
    port map (
            O => \N__1435\,
            I => \N__1431\
        );

    \I__237\ : InMux
    port map (
            O => \N__1434\,
            I => \N__1428\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__1431\,
            I => \N__1425\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1428\,
            I => \cntDivZ0Z_20\
        );

    \I__234\ : Odrv4
    port map (
            O => \N__1425\,
            I => \cntDivZ0Z_20\
        );

    \I__233\ : CascadeMux
    port map (
            O => \N__1420\,
            I => \N__1417\
        );

    \I__232\ : InMux
    port map (
            O => \N__1417\,
            I => \N__1413\
        );

    \I__231\ : InMux
    port map (
            O => \N__1416\,
            I => \N__1410\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__1413\,
            I => \N__1407\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__1410\,
            I => \cntDivZ0Z_21\
        );

    \I__228\ : Odrv4
    port map (
            O => \N__1407\,
            I => \cntDivZ0Z_21\
        );

    \I__227\ : CascadeMux
    port map (
            O => \N__1402\,
            I => \N__1399\
        );

    \I__226\ : InMux
    port map (
            O => \N__1399\,
            I => \N__1395\
        );

    \I__225\ : InMux
    port map (
            O => \N__1398\,
            I => \N__1392\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1395\,
            I => \N__1389\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1392\,
            I => \cntDivZ0Z_22\
        );

    \I__222\ : Odrv4
    port map (
            O => \N__1389\,
            I => \cntDivZ0Z_22\
        );

    \I__221\ : CascadeMux
    port map (
            O => \N__1384\,
            I => \N__1381\
        );

    \I__220\ : InMux
    port map (
            O => \N__1381\,
            I => \N__1377\
        );

    \I__219\ : InMux
    port map (
            O => \N__1380\,
            I => \N__1374\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1377\,
            I => \N__1371\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__1374\,
            I => \cntDivZ0Z_23\
        );

    \I__216\ : Odrv4
    port map (
            O => \N__1371\,
            I => \cntDivZ0Z_23\
        );

    \I__215\ : InMux
    port map (
            O => \N__1366\,
            I => \N__1362\
        );

    \I__214\ : InMux
    port map (
            O => \N__1365\,
            I => \N__1359\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1362\,
            I => \N__1356\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1359\,
            I => \cntDivZ0Z_24\
        );

    \I__211\ : Odrv4
    port map (
            O => \N__1356\,
            I => \cntDivZ0Z_24\
        );

    \I__210\ : CascadeMux
    port map (
            O => \N__1351\,
            I => \N__1348\
        );

    \I__209\ : InMux
    port map (
            O => \N__1348\,
            I => \N__1344\
        );

    \I__208\ : InMux
    port map (
            O => \N__1347\,
            I => \N__1341\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1344\,
            I => \N__1338\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__1341\,
            I => \cntDivZ0Z_8\
        );

    \I__205\ : Odrv4
    port map (
            O => \N__1338\,
            I => \cntDivZ0Z_8\
        );

    \I__204\ : CascadeMux
    port map (
            O => \N__1333\,
            I => \N__1330\
        );

    \I__203\ : InMux
    port map (
            O => \N__1330\,
            I => \N__1326\
        );

    \I__202\ : InMux
    port map (
            O => \N__1329\,
            I => \N__1323\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1326\,
            I => \N__1320\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__1323\,
            I => \cntDivZ0Z_9\
        );

    \I__199\ : Odrv12
    port map (
            O => \N__1320\,
            I => \cntDivZ0Z_9\
        );

    \I__198\ : CascadeMux
    port map (
            O => \N__1315\,
            I => \N__1312\
        );

    \I__197\ : InMux
    port map (
            O => \N__1312\,
            I => \N__1308\
        );

    \I__196\ : InMux
    port map (
            O => \N__1311\,
            I => \N__1305\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1308\,
            I => \N__1302\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1305\,
            I => \cntDivZ0Z_10\
        );

    \I__193\ : Odrv12
    port map (
            O => \N__1302\,
            I => \cntDivZ0Z_10\
        );

    \I__192\ : CascadeMux
    port map (
            O => \N__1297\,
            I => \N__1294\
        );

    \I__191\ : InMux
    port map (
            O => \N__1294\,
            I => \N__1290\
        );

    \I__190\ : InMux
    port map (
            O => \N__1293\,
            I => \N__1287\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1290\,
            I => \N__1284\
        );

    \I__188\ : LocalMux
    port map (
            O => \N__1287\,
            I => \cntDivZ0Z_11\
        );

    \I__187\ : Odrv4
    port map (
            O => \N__1284\,
            I => \cntDivZ0Z_11\
        );

    \I__186\ : InMux
    port map (
            O => \N__1279\,
            I => \N__1275\
        );

    \I__185\ : InMux
    port map (
            O => \N__1278\,
            I => \N__1272\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1275\,
            I => \N__1269\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1272\,
            I => \cntDivZ0Z_12\
        );

    \I__182\ : Odrv4
    port map (
            O => \N__1269\,
            I => \cntDivZ0Z_12\
        );

    \I__181\ : CascadeMux
    port map (
            O => \N__1264\,
            I => \N__1261\
        );

    \I__180\ : InMux
    port map (
            O => \N__1261\,
            I => \N__1257\
        );

    \I__179\ : InMux
    port map (
            O => \N__1260\,
            I => \N__1254\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1257\,
            I => \N__1251\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1254\,
            I => \cntDivZ0Z_13\
        );

    \I__176\ : Odrv4
    port map (
            O => \N__1251\,
            I => \cntDivZ0Z_13\
        );

    \I__175\ : CascadeMux
    port map (
            O => \N__1246\,
            I => \N__1243\
        );

    \I__174\ : InMux
    port map (
            O => \N__1243\,
            I => \N__1239\
        );

    \I__173\ : InMux
    port map (
            O => \N__1242\,
            I => \N__1236\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1239\,
            I => \N__1233\
        );

    \I__171\ : LocalMux
    port map (
            O => \N__1236\,
            I => \cntDivZ0Z_14\
        );

    \I__170\ : Odrv4
    port map (
            O => \N__1233\,
            I => \cntDivZ0Z_14\
        );

    \I__169\ : CascadeMux
    port map (
            O => \N__1228\,
            I => \N__1225\
        );

    \I__168\ : InMux
    port map (
            O => \N__1225\,
            I => \N__1221\
        );

    \I__167\ : InMux
    port map (
            O => \N__1224\,
            I => \N__1218\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1221\,
            I => \N__1215\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__1218\,
            I => \cntDivZ0Z_15\
        );

    \I__164\ : Odrv4
    port map (
            O => \N__1215\,
            I => \cntDivZ0Z_15\
        );

    \I__163\ : InMux
    port map (
            O => \N__1210\,
            I => un2_cntdiv_cry_22
        );

    \I__162\ : InMux
    port map (
            O => \N__1207\,
            I => un2_cntdiv_cry_23
        );

    \I__161\ : CascadeMux
    port map (
            O => \N__1204\,
            I => \N__1201\
        );

    \I__160\ : InMux
    port map (
            O => \N__1201\,
            I => \N__1196\
        );

    \I__159\ : InMux
    port map (
            O => \N__1200\,
            I => \N__1190\
        );

    \I__158\ : InMux
    port map (
            O => \N__1199\,
            I => \N__1190\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__1196\,
            I => \N__1187\
        );

    \I__156\ : InMux
    port map (
            O => \N__1195\,
            I => \N__1184\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__1190\,
            I => \cntDivZ0Z_0\
        );

    \I__154\ : Odrv4
    port map (
            O => \N__1187\,
            I => \cntDivZ0Z_0\
        );

    \I__153\ : LocalMux
    port map (
            O => \N__1184\,
            I => \cntDivZ0Z_0\
        );

    \I__152\ : InMux
    port map (
            O => \N__1177\,
            I => \N__1172\
        );

    \I__151\ : CascadeMux
    port map (
            O => \N__1176\,
            I => \N__1169\
        );

    \I__150\ : InMux
    port map (
            O => \N__1175\,
            I => \N__1166\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__1172\,
            I => \N__1163\
        );

    \I__148\ : InMux
    port map (
            O => \N__1169\,
            I => \N__1160\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1166\,
            I => \cntDivZ0Z_1\
        );

    \I__146\ : Odrv4
    port map (
            O => \N__1163\,
            I => \cntDivZ0Z_1\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1160\,
            I => \cntDivZ0Z_1\
        );

    \I__144\ : CascadeMux
    port map (
            O => \N__1153\,
            I => \N__1150\
        );

    \I__143\ : InMux
    port map (
            O => \N__1150\,
            I => \N__1146\
        );

    \I__142\ : InMux
    port map (
            O => \N__1149\,
            I => \N__1143\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1146\,
            I => \N__1140\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1143\,
            I => \cntDivZ0Z_2\
        );

    \I__139\ : Odrv12
    port map (
            O => \N__1140\,
            I => \cntDivZ0Z_2\
        );

    \I__138\ : InMux
    port map (
            O => \N__1135\,
            I => \N__1131\
        );

    \I__137\ : InMux
    port map (
            O => \N__1134\,
            I => \N__1128\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__1131\,
            I => \N__1125\
        );

    \I__135\ : LocalMux
    port map (
            O => \N__1128\,
            I => \cntDivZ0Z_3\
        );

    \I__134\ : Odrv4
    port map (
            O => \N__1125\,
            I => \cntDivZ0Z_3\
        );

    \I__133\ : CascadeMux
    port map (
            O => \N__1120\,
            I => \N__1117\
        );

    \I__132\ : InMux
    port map (
            O => \N__1117\,
            I => \N__1113\
        );

    \I__131\ : InMux
    port map (
            O => \N__1116\,
            I => \N__1110\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__1113\,
            I => \N__1107\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1110\,
            I => \cntDivZ0Z_4\
        );

    \I__128\ : Odrv4
    port map (
            O => \N__1107\,
            I => \cntDivZ0Z_4\
        );

    \I__127\ : CascadeMux
    port map (
            O => \N__1102\,
            I => \N__1099\
        );

    \I__126\ : InMux
    port map (
            O => \N__1099\,
            I => \N__1095\
        );

    \I__125\ : InMux
    port map (
            O => \N__1098\,
            I => \N__1092\
        );

    \I__124\ : LocalMux
    port map (
            O => \N__1095\,
            I => \N__1089\
        );

    \I__123\ : LocalMux
    port map (
            O => \N__1092\,
            I => \cntDivZ0Z_5\
        );

    \I__122\ : Odrv4
    port map (
            O => \N__1089\,
            I => \cntDivZ0Z_5\
        );

    \I__121\ : CascadeMux
    port map (
            O => \N__1084\,
            I => \N__1081\
        );

    \I__120\ : InMux
    port map (
            O => \N__1081\,
            I => \N__1077\
        );

    \I__119\ : InMux
    port map (
            O => \N__1080\,
            I => \N__1074\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__1077\,
            I => \N__1071\
        );

    \I__117\ : LocalMux
    port map (
            O => \N__1074\,
            I => \cntDivZ0Z_6\
        );

    \I__116\ : Odrv4
    port map (
            O => \N__1071\,
            I => \cntDivZ0Z_6\
        );

    \I__115\ : CascadeMux
    port map (
            O => \N__1066\,
            I => \N__1063\
        );

    \I__114\ : InMux
    port map (
            O => \N__1063\,
            I => \N__1059\
        );

    \I__113\ : InMux
    port map (
            O => \N__1062\,
            I => \N__1056\
        );

    \I__112\ : LocalMux
    port map (
            O => \N__1059\,
            I => \N__1053\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__1056\,
            I => \cntDivZ0Z_7\
        );

    \I__110\ : Odrv4
    port map (
            O => \N__1053\,
            I => \cntDivZ0Z_7\
        );

    \I__109\ : InMux
    port map (
            O => \N__1048\,
            I => un2_cntdiv_cry_13
        );

    \I__108\ : InMux
    port map (
            O => \N__1045\,
            I => un2_cntdiv_cry_14
        );

    \I__107\ : InMux
    port map (
            O => \N__1042\,
            I => un2_cntdiv_cry_15
        );

    \I__106\ : InMux
    port map (
            O => \N__1039\,
            I => \bfn_22_19_0_\
        );

    \I__105\ : InMux
    port map (
            O => \N__1036\,
            I => un2_cntdiv_cry_17
        );

    \I__104\ : InMux
    port map (
            O => \N__1033\,
            I => un2_cntdiv_cry_18
        );

    \I__103\ : InMux
    port map (
            O => \N__1030\,
            I => un2_cntdiv_cry_19
        );

    \I__102\ : InMux
    port map (
            O => \N__1027\,
            I => un2_cntdiv_cry_20
        );

    \I__101\ : InMux
    port map (
            O => \N__1024\,
            I => un2_cntdiv_cry_21
        );

    \I__100\ : InMux
    port map (
            O => \N__1021\,
            I => un2_cntdiv_cry_4
        );

    \I__99\ : InMux
    port map (
            O => \N__1018\,
            I => un2_cntdiv_cry_5
        );

    \I__98\ : InMux
    port map (
            O => \N__1015\,
            I => un2_cntdiv_cry_6
        );

    \I__97\ : InMux
    port map (
            O => \N__1012\,
            I => un2_cntdiv_cry_7
        );

    \I__96\ : InMux
    port map (
            O => \N__1009\,
            I => \bfn_22_18_0_\
        );

    \I__95\ : InMux
    port map (
            O => \N__1006\,
            I => un2_cntdiv_cry_9
        );

    \I__94\ : InMux
    port map (
            O => \N__1003\,
            I => un2_cntdiv_cry_10
        );

    \I__93\ : InMux
    port map (
            O => \N__1000\,
            I => un2_cntdiv_cry_11
        );

    \I__92\ : InMux
    port map (
            O => \N__997\,
            I => un2_cntdiv_cry_12
        );

    \I__91\ : InMux
    port map (
            O => \N__994\,
            I => un2_cntdiv_cry_1
        );

    \I__90\ : InMux
    port map (
            O => \N__991\,
            I => un2_cntdiv_cry_2
        );

    \I__89\ : InMux
    port map (
            O => \N__988\,
            I => un2_cntdiv_cry_3
        );

    \IN_MUX_bfv_22_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_17_0_\
        );

    \IN_MUX_bfv_22_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_cntdiv_cry_8,
            carryinitout => \bfn_22_18_0_\
        );

    \IN_MUX_bfv_22_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_cntdiv_cry_16,
            carryinitout => \bfn_22_19_0_\
        );

    \IN_MUX_bfv_22_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_20_0_\
        );

    \IN_MUX_bfv_22_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_cntdiv_1_cry_8,
            carryinitout => \bfn_22_21_0_\
        );

    \IN_MUX_bfv_22_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_cntdiv_1_cry_16,
            carryinitout => \bfn_22_22_0_\
        );

    \IN_MUX_bfv_22_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_cntdiv_1_cry_24,
            carryinitout => \bfn_22_23_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \cntDiv_1_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1199\,
            in2 => \_gnd_net_\,
            in3 => \N__1175\,
            lcout => \cntDivZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_0_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cntDivZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_cry_1_c_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1177\,
            in2 => \N__1204\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_17_0_\,
            carryout => un2_cntdiv_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_2_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1149\,
            in2 => \_gnd_net_\,
            in3 => \N__994\,
            lcout => \cntDivZ0Z_2\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_1,
            carryout => un2_cntdiv_cry_2,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_3_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1134\,
            in2 => \_gnd_net_\,
            in3 => \N__991\,
            lcout => \cntDivZ0Z_3\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_2,
            carryout => un2_cntdiv_cry_3,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_4_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1116\,
            in2 => \_gnd_net_\,
            in3 => \N__988\,
            lcout => \cntDivZ0Z_4\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_3,
            carryout => un2_cntdiv_cry_4,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_5_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1098\,
            in2 => \_gnd_net_\,
            in3 => \N__1021\,
            lcout => \cntDivZ0Z_5\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_4,
            carryout => un2_cntdiv_cry_5,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_6_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1080\,
            in2 => \_gnd_net_\,
            in3 => \N__1018\,
            lcout => \cntDivZ0Z_6\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_5,
            carryout => un2_cntdiv_cry_6,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_7_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1062\,
            in2 => \_gnd_net_\,
            in3 => \N__1015\,
            lcout => \cntDivZ0Z_7\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_6,
            carryout => un2_cntdiv_cry_7,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_8_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1347\,
            in2 => \_gnd_net_\,
            in3 => \N__1012\,
            lcout => \cntDivZ0Z_8\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_7,
            carryout => un2_cntdiv_cry_8,
            clk => \N__1578\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_9_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1329\,
            in2 => \_gnd_net_\,
            in3 => \N__1009\,
            lcout => \cntDivZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_22_18_0_\,
            carryout => un2_cntdiv_cry_9,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_10_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1311\,
            in2 => \_gnd_net_\,
            in3 => \N__1006\,
            lcout => \cntDivZ0Z_10\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_9,
            carryout => un2_cntdiv_cry_10,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_11_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1293\,
            in2 => \_gnd_net_\,
            in3 => \N__1003\,
            lcout => \cntDivZ0Z_11\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_10,
            carryout => un2_cntdiv_cry_11,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_12_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1278\,
            in2 => \_gnd_net_\,
            in3 => \N__1000\,
            lcout => \cntDivZ0Z_12\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_11,
            carryout => un2_cntdiv_cry_12,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_13_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1260\,
            in2 => \_gnd_net_\,
            in3 => \N__997\,
            lcout => \cntDivZ0Z_13\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_12,
            carryout => un2_cntdiv_cry_13,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_14_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1242\,
            in2 => \_gnd_net_\,
            in3 => \N__1048\,
            lcout => \cntDivZ0Z_14\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_13,
            carryout => un2_cntdiv_cry_14,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_15_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1224\,
            in2 => \_gnd_net_\,
            in3 => \N__1045\,
            lcout => \cntDivZ0Z_15\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_14,
            carryout => un2_cntdiv_cry_15,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_16_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1506\,
            in2 => \_gnd_net_\,
            in3 => \N__1042\,
            lcout => \cntDivZ0Z_16\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_15,
            carryout => un2_cntdiv_cry_16,
            clk => \N__1579\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_17_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1488\,
            in2 => \_gnd_net_\,
            in3 => \N__1039\,
            lcout => \cntDivZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_22_19_0_\,
            carryout => un2_cntdiv_cry_17,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_18_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1470\,
            in2 => \_gnd_net_\,
            in3 => \N__1036\,
            lcout => \cntDivZ0Z_18\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_17,
            carryout => un2_cntdiv_cry_18,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_19_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1452\,
            in2 => \_gnd_net_\,
            in3 => \N__1033\,
            lcout => \cntDivZ0Z_19\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_18,
            carryout => un2_cntdiv_cry_19,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_20_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1434\,
            in2 => \_gnd_net_\,
            in3 => \N__1030\,
            lcout => \cntDivZ0Z_20\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_19,
            carryout => un2_cntdiv_cry_20,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_21_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1416\,
            in2 => \_gnd_net_\,
            in3 => \N__1027\,
            lcout => \cntDivZ0Z_21\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_20,
            carryout => un2_cntdiv_cry_21,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_22_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1398\,
            in2 => \_gnd_net_\,
            in3 => \N__1024\,
            lcout => \cntDivZ0Z_22\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_21,
            carryout => un2_cntdiv_cry_22,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_23_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1380\,
            in2 => \_gnd_net_\,
            in3 => \N__1210\,
            lcout => \cntDivZ0Z_23\,
            ltout => OPEN,
            carryin => un2_cntdiv_cry_22,
            carryout => un2_cntdiv_cry_23,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_24_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1365\,
            in2 => \_gnd_net_\,
            in3 => \N__1207\,
            lcout => \cntDivZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1581\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_1_c_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1195\,
            in2 => \N__1176\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_20_0_\,
            carryout => un2_cntdiv_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_2_c_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1153\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_1,
            carryout => un2_cntdiv_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_3_c_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1135\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_2,
            carryout => un2_cntdiv_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_4_c_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_3,
            carryout => un2_cntdiv_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_5_c_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1102\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_4,
            carryout => un2_cntdiv_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_6_c_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1084\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_5,
            carryout => un2_cntdiv_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_7_c_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1066\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_6,
            carryout => un2_cntdiv_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_8_c_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1351\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_7,
            carryout => un2_cntdiv_1_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_9_c_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1333\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_21_0_\,
            carryout => un2_cntdiv_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_10_c_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1315\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_9,
            carryout => un2_cntdiv_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_11_c_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1297\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_10,
            carryout => un2_cntdiv_1_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_12_c_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1279\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_11,
            carryout => un2_cntdiv_1_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_13_c_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1264\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_12,
            carryout => un2_cntdiv_1_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_14_c_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1246\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_13,
            carryout => un2_cntdiv_1_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_15_c_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1228\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_14,
            carryout => un2_cntdiv_1_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_16_c_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1510\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_15,
            carryout => un2_cntdiv_1_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_17_c_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1492\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_22_22_0_\,
            carryout => un2_cntdiv_1_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_18_c_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1474\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_17,
            carryout => un2_cntdiv_1_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_19_c_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1456\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_18,
            carryout => un2_cntdiv_1_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_20_c_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1438\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_19,
            carryout => un2_cntdiv_1_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_21_c_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1420\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_20,
            carryout => un2_cntdiv_1_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_22_c_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1402\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_21,
            carryout => un2_cntdiv_1_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_23_c_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1384\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_22,
            carryout => un2_cntdiv_1_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_24_c_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1366\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un2_cntdiv_1_cry_23,
            carryout => un2_cntdiv_1_cry_24,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_cntdiv_1_cry_24_c_RNI73PB_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1596\,
            in2 => \_gnd_net_\,
            in3 => \N__1612\,
            lcout => \un2_cntdiv_1_cry_24_c_RNI73PBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter1.Pre_Q_1_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__1811\,
            in1 => \N__1879\,
            in2 => \_gnd_net_\,
            in3 => \N__1678\,
            lcout => value_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1582\,
            ce => \N__1551\,
            sr => \_gnd_net_\
        );

    \cntDiv_RNIETOH_25_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1597\,
            in2 => \_gnd_net_\,
            in3 => \N__1608\,
            lcout => \cntDiv_RNIETOHZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntDiv_25_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1609\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cntDiv_i_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1584\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter1.Pre_Q_3_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000010"
        )
    port map (
            in0 => \N__1812\,
            in1 => \N__1880\,
            in2 => \N__1691\,
            in3 => \N__1741\,
            lcout => value_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1583\,
            ce => \N__1555\,
            sr => \_gnd_net_\
        );

    \counter1.Pre_Q_2_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__1673\,
            in1 => \N__1814\,
            in2 => \N__1898\,
            in3 => \N__1740\,
            lcout => value_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1585\,
            ce => \N__1550\,
            sr => \_gnd_net_\
        );

    \counter1.Pre_Q_0_LC_24_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__1813\,
            in1 => \N__1881\,
            in2 => \N__1748\,
            in3 => \N__1674\,
            lcout => value_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__1585\,
            ce => \N__1550\,
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m6_LC_32_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101100110"
        )
    port map (
            in0 => \N__1783\,
            in1 => \N__1830\,
            in2 => \N__1714\,
            in3 => \N__1903\,
            lcout => \Y_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m15_LC_32_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100100100"
        )
    port map (
            in0 => \N__1781\,
            in1 => \N__1828\,
            in2 => \N__1713\,
            in3 => \N__1902\,
            lcout => \Y_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m2_LC_32_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__1829\,
            in1 => \N__1782\,
            in2 => \_gnd_net_\,
            in3 => \N__1904\,
            lcout => \Y_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m11_LC_32_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001000110"
        )
    port map (
            in0 => \N__1827\,
            in1 => \N__1780\,
            in2 => \N__1908\,
            in3 => \N__1706\,
            lcout => \Y_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m19_LC_32_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100111000"
        )
    port map (
            in0 => \N__1695\,
            in1 => \N__1768\,
            in2 => \N__1852\,
            in3 => \N__1921\,
            lcout => \Y_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m18_LC_32_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100010110"
        )
    port map (
            in0 => \N__1920\,
            in1 => \N__1847\,
            in2 => \N__1779\,
            in3 => \N__1694\,
            lcout => \Y_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m13_LC_32_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010000"
        )
    port map (
            in0 => \N__1692\,
            in1 => \N__1761\,
            in2 => \N__1851\,
            in3 => \N__1918\,
            lcout => \Y_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \display.S_1_7_0__m16_LC_32_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110100"
        )
    port map (
            in0 => \N__1919\,
            in1 => \N__1846\,
            in2 => \N__1778\,
            in3 => \N__1693\,
            lcout => \Y_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_32_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
